VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO mem_64_32_gf180
  FOREIGN mem_64_32_gf180 0 0 ;
  CLASS BLOCK ;
  SIZE 1020 BY 620 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  992.26 14.546 996.74 257.614 ;
        RECT  11.48 347.186 13.72 590.254 ;
        RECT  992.26 347.186 996.74 590.254 ;
        RECT  11.48 14.546 13.72 257.614 ;
        RECT  976.08 14.546 980.56 610.414 ;
        RECT  931.28 14.546 935.76 610.414 ;
        RECT  886.48 14.546 890.96 610.414 ;
        RECT  841.68 14.546 846.16 610.414 ;
        RECT  796.88 14.546 801.36 610.414 ;
        RECT  752.08 14.546 756.56 610.414 ;
        RECT  707.28 14.546 711.76 610.414 ;
        RECT  662.48 14.546 666.96 610.414 ;
        RECT  617.68 14.546 622.16 610.414 ;
        RECT  572.88 14.546 577.36 610.414 ;
        RECT  528.08 14.546 532.56 610.414 ;
        RECT  483.28 14.546 487.76 610.414 ;
        RECT  438.48 14.546 442.96 610.414 ;
        RECT  393.68 14.546 398.16 610.414 ;
        RECT  348.88 14.546 353.36 610.414 ;
        RECT  304.08 14.546 308.56 610.414 ;
        RECT  259.28 14.546 263.76 610.414 ;
        RECT  214.48 14.546 218.96 610.414 ;
        RECT  169.68 14.546 174.16 610.414 ;
        RECT  124.88 14.546 129.36 610.414 ;
        RECT  80.08 14.546 84.56 610.414 ;
        RECT  35.28 14.546 39.76 610.414 ;
      LAYER Metal1 ;
        RECT  985.04 579.15 1009.68 580.05 ;
        RECT  985.04 569.07 1009.68 569.97 ;
        RECT  985.04 558.99 1009.68 559.89 ;
        RECT  985.04 548.91 1009.68 549.81 ;
        RECT  985.04 538.83 1009.68 539.73 ;
        RECT  985.04 528.75 1009.68 529.65 ;
        RECT  985.04 518.67 1009.68 519.57 ;
        RECT  985.04 508.59 1009.68 509.49 ;
        RECT  985.04 498.51 1009.68 499.41 ;
        RECT  985.04 488.43 1009.68 489.33 ;
        RECT  985.04 478.35 1009.68 479.25 ;
        RECT  985.04 468.27 1009.68 469.17 ;
        RECT  985.04 458.19 1009.68 459.09 ;
        RECT  985.04 448.11 1009.68 449.01 ;
        RECT  985.04 438.03 1009.68 438.93 ;
        RECT  985.04 427.95 1009.68 428.85 ;
        RECT  985.04 417.87 1009.68 418.77 ;
        RECT  985.04 407.79 1009.68 408.69 ;
        RECT  985.04 397.71 1009.68 398.61 ;
        RECT  985.04 387.63 1009.68 388.53 ;
        RECT  985.04 377.55 1009.68 378.45 ;
        RECT  985.04 367.47 1009.68 368.37 ;
        RECT  985.04 357.39 1009.68 358.29 ;
        RECT  985.04 246.51 1009.68 247.41 ;
        RECT  985.04 236.43 1009.68 237.33 ;
        RECT  985.04 226.35 1009.68 227.25 ;
        RECT  985.04 216.27 1009.68 217.17 ;
        RECT  985.04 206.19 1009.68 207.09 ;
        RECT  985.04 196.11 1009.68 197.01 ;
        RECT  985.04 186.03 1009.68 186.93 ;
        RECT  985.04 175.95 1009.68 176.85 ;
        RECT  985.04 165.87 1009.68 166.77 ;
        RECT  985.04 155.79 1009.68 156.69 ;
        RECT  985.04 145.71 1009.68 146.61 ;
        RECT  985.04 135.63 1009.68 136.53 ;
        RECT  985.04 125.55 1009.68 126.45 ;
        RECT  985.04 115.47 1009.68 116.37 ;
        RECT  985.04 105.39 1009.68 106.29 ;
        RECT  985.04 95.31 1009.68 96.21 ;
        RECT  985.04 85.23 1009.68 86.13 ;
        RECT  985.04 75.15 1009.68 76.05 ;
        RECT  985.04 65.07 1009.68 65.97 ;
        RECT  985.04 54.99 1009.68 55.89 ;
        RECT  985.04 44.91 1009.68 45.81 ;
        RECT  985.04 34.83 1009.68 35.73 ;
        RECT  985.04 24.75 1009.68 25.65 ;
        RECT  454.16 579.15 548.8 580.05 ;
        RECT  454.16 569.07 548.8 569.97 ;
        RECT  454.16 558.99 548.8 559.89 ;
        RECT  454.16 548.91 548.8 549.81 ;
        RECT  454.16 538.83 548.8 539.73 ;
        RECT  454.16 528.75 548.8 529.65 ;
        RECT  454.16 518.67 548.8 519.57 ;
        RECT  454.16 508.59 548.8 509.49 ;
        RECT  454.16 498.51 548.8 499.41 ;
        RECT  454.16 488.43 548.8 489.33 ;
        RECT  454.16 478.35 548.8 479.25 ;
        RECT  454.16 468.27 548.8 469.17 ;
        RECT  454.16 458.19 548.8 459.09 ;
        RECT  454.16 448.11 548.8 449.01 ;
        RECT  454.16 438.03 548.8 438.93 ;
        RECT  454.16 427.95 548.8 428.85 ;
        RECT  454.16 417.87 548.8 418.77 ;
        RECT  454.16 407.79 548.8 408.69 ;
        RECT  454.16 397.71 548.8 398.61 ;
        RECT  454.16 387.63 548.8 388.53 ;
        RECT  454.16 377.55 548.8 378.45 ;
        RECT  454.16 367.47 548.8 368.37 ;
        RECT  454.16 357.39 548.8 358.29 ;
        RECT  454.16 246.51 548.8 247.41 ;
        RECT  454.16 236.43 548.8 237.33 ;
        RECT  454.16 226.35 548.8 227.25 ;
        RECT  454.16 216.27 548.8 217.17 ;
        RECT  454.16 206.19 548.8 207.09 ;
        RECT  454.16 196.11 548.8 197.01 ;
        RECT  454.16 186.03 548.8 186.93 ;
        RECT  454.16 175.95 548.8 176.85 ;
        RECT  454.16 165.87 548.8 166.77 ;
        RECT  454.16 155.79 548.8 156.69 ;
        RECT  454.16 145.71 548.8 146.61 ;
        RECT  454.16 135.63 548.8 136.53 ;
        RECT  454.16 125.55 548.8 126.45 ;
        RECT  454.16 115.47 548.8 116.37 ;
        RECT  454.16 105.39 548.8 106.29 ;
        RECT  454.16 95.31 548.8 96.21 ;
        RECT  454.16 85.23 548.8 86.13 ;
        RECT  454.16 75.15 548.8 76.05 ;
        RECT  454.16 65.07 548.8 65.97 ;
        RECT  454.16 54.99 548.8 55.89 ;
        RECT  454.16 44.91 548.8 45.81 ;
        RECT  454.16 34.83 548.8 35.73 ;
        RECT  454.16 24.75 548.8 25.65 ;
        RECT  10.08 609.39 1009.68 610.29 ;
        RECT  10.08 599.31 1009.68 600.21 ;
        RECT  10.08 589.23 1009.68 590.13 ;
        RECT  10.08 579.15 17.92 580.05 ;
        RECT  10.08 569.07 17.92 569.97 ;
        RECT  10.08 558.99 17.92 559.89 ;
        RECT  10.08 548.91 17.92 549.81 ;
        RECT  10.08 538.83 17.92 539.73 ;
        RECT  10.08 528.75 17.92 529.65 ;
        RECT  10.08 518.67 17.92 519.57 ;
        RECT  10.08 508.59 17.92 509.49 ;
        RECT  10.08 498.51 17.92 499.41 ;
        RECT  10.08 488.43 17.92 489.33 ;
        RECT  10.08 478.35 17.92 479.25 ;
        RECT  10.08 468.27 17.92 469.17 ;
        RECT  10.08 458.19 17.92 459.09 ;
        RECT  10.08 448.11 17.92 449.01 ;
        RECT  10.08 438.03 17.92 438.93 ;
        RECT  10.08 427.95 17.92 428.85 ;
        RECT  10.08 417.87 17.92 418.77 ;
        RECT  10.08 407.79 17.92 408.69 ;
        RECT  10.08 397.71 17.92 398.61 ;
        RECT  10.08 387.63 17.92 388.53 ;
        RECT  10.08 377.55 17.92 378.45 ;
        RECT  10.08 367.47 17.92 368.37 ;
        RECT  10.08 357.39 17.92 358.29 ;
        RECT  10.08 347.31 1009.68 348.21 ;
        RECT  10.08 337.23 1009.68 338.13 ;
        RECT  10.08 327.15 1009.68 328.05 ;
        RECT  10.08 317.07 1009.68 317.97 ;
        RECT  10.08 306.99 1009.68 307.89 ;
        RECT  10.08 296.91 1009.68 297.81 ;
        RECT  10.08 286.83 1009.68 287.73 ;
        RECT  10.08 276.75 1009.68 277.65 ;
        RECT  10.08 266.67 1009.68 267.57 ;
        RECT  10.08 256.59 1009.68 257.49 ;
        RECT  10.08 246.51 17.92 247.41 ;
        RECT  10.08 236.43 17.92 237.33 ;
        RECT  10.08 226.35 17.92 227.25 ;
        RECT  10.08 216.27 17.92 217.17 ;
        RECT  10.08 206.19 17.92 207.09 ;
        RECT  10.08 196.11 17.92 197.01 ;
        RECT  10.08 186.03 17.92 186.93 ;
        RECT  10.08 175.95 17.92 176.85 ;
        RECT  10.08 165.87 17.92 166.77 ;
        RECT  10.08 155.79 17.92 156.69 ;
        RECT  10.08 145.71 17.92 146.61 ;
        RECT  10.08 135.63 17.92 136.53 ;
        RECT  10.08 125.55 17.92 126.45 ;
        RECT  10.08 115.47 17.92 116.37 ;
        RECT  10.08 105.39 17.92 106.29 ;
        RECT  10.08 95.31 17.92 96.21 ;
        RECT  10.08 85.23 17.92 86.13 ;
        RECT  10.08 75.15 17.92 76.05 ;
        RECT  10.08 65.07 17.92 65.97 ;
        RECT  10.08 54.99 17.92 55.89 ;
        RECT  10.08 44.91 17.92 45.81 ;
        RECT  10.08 34.83 17.92 35.73 ;
        RECT  10.08 24.75 17.92 25.65 ;
        RECT  10.08 14.67 1009.68 15.57 ;
      VIA 994.756 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 589.106 995.63 590.254 ;
      VIA 994.816 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 579.026 995.63 580.174 ;
      VIA 994.816 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 568.946 995.63 570.094 ;
      VIA 994.816 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 558.866 995.63 560.014 ;
      VIA 994.816 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 548.786 995.63 549.934 ;
      VIA 994.816 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 538.706 995.63 539.854 ;
      VIA 994.816 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 528.626 995.63 529.774 ;
      VIA 994.816 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 518.546 995.63 519.694 ;
      VIA 994.816 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 508.466 995.63 509.614 ;
      VIA 994.816 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 498.386 995.63 499.534 ;
      VIA 994.816 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 488.306 995.63 489.454 ;
      VIA 994.816 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 478.226 995.63 479.374 ;
      VIA 994.816 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 468.146 995.63 469.294 ;
      VIA 994.816 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 458.066 995.63 459.214 ;
      VIA 994.816 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 447.986 995.63 449.134 ;
      VIA 994.816 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 437.906 995.63 439.054 ;
      VIA 994.816 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 427.826 995.63 428.974 ;
      VIA 994.816 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 417.746 995.63 418.894 ;
      VIA 994.816 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 407.666 995.63 408.814 ;
      VIA 994.816 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 397.586 995.63 398.734 ;
      VIA 994.816 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 387.506 995.63 388.654 ;
      VIA 994.816 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 377.426 995.63 378.574 ;
      VIA 994.816 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 367.346 995.63 368.494 ;
      VIA 994.816 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 357.266 995.63 358.414 ;
      VIA 994.816 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 347.186 995.63 348.334 ;
      VIA 994.816 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 256.466 995.63 257.614 ;
      VIA 994.816 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 246.386 995.63 247.534 ;
      VIA 994.816 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 236.306 995.63 237.454 ;
      VIA 994.816 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 226.226 995.63 227.374 ;
      VIA 994.816 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 216.146 995.63 217.294 ;
      VIA 994.816 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 206.066 995.63 207.214 ;
      VIA 994.816 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 195.986 995.63 197.134 ;
      VIA 994.816 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 185.906 995.63 187.054 ;
      VIA 994.816 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 175.826 995.63 176.974 ;
      VIA 994.816 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 165.746 995.63 166.894 ;
      VIA 994.816 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 155.666 995.63 156.814 ;
      VIA 994.816 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 145.586 995.63 146.734 ;
      VIA 994.816 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 135.506 995.63 136.654 ;
      VIA 994.816 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 125.426 995.63 126.574 ;
      VIA 994.816 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 115.346 995.63 116.494 ;
      VIA 994.816 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 105.266 995.63 106.414 ;
      VIA 994.816 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 95.186 995.63 96.334 ;
      VIA 994.816 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 85.106 995.63 86.254 ;
      VIA 994.816 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 75.026 995.63 76.174 ;
      VIA 994.816 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 64.946 995.63 66.094 ;
      VIA 994.816 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 54.866 995.63 56.014 ;
      VIA 994.816 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 44.786 995.63 45.934 ;
      VIA 994.816 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 34.706 995.63 35.854 ;
      VIA 994.816 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 24.626 995.63 25.774 ;
      VIA 994.816 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 994.756 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.756 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.628 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.5 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.372 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 994.244 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  993.49 14.546 995.63 15.694 ;
      VIA 994.816 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.816 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.688 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.432 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.304 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 994.56 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 609.266 979.39 610.414 ;
      VIA 978.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 599.186 979.39 600.334 ;
      VIA 978.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 589.106 979.39 590.254 ;
      VIA 978.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 347.186 979.39 348.334 ;
      VIA 978.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 337.106 979.39 338.254 ;
      VIA 978.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 327.026 979.39 328.174 ;
      VIA 978.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 316.946 979.39 318.094 ;
      VIA 978.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 306.866 979.39 308.014 ;
      VIA 978.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 296.786 979.39 297.934 ;
      VIA 978.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 286.706 979.39 287.854 ;
      VIA 978.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 276.626 979.39 277.774 ;
      VIA 978.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 266.546 979.39 267.694 ;
      VIA 978.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 256.466 979.39 257.614 ;
      VIA 978.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 978.556 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.556 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.428 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.3 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.172 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 978.044 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  977.25 14.546 979.39 15.694 ;
      VIA 978.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 978.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 609.266 934.59 610.414 ;
      VIA 933.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 599.186 934.59 600.334 ;
      VIA 933.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 589.106 934.59 590.254 ;
      VIA 933.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 347.186 934.59 348.334 ;
      VIA 933.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 337.106 934.59 338.254 ;
      VIA 933.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 327.026 934.59 328.174 ;
      VIA 933.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 316.946 934.59 318.094 ;
      VIA 933.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 306.866 934.59 308.014 ;
      VIA 933.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 296.786 934.59 297.934 ;
      VIA 933.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 286.706 934.59 287.854 ;
      VIA 933.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 276.626 934.59 277.774 ;
      VIA 933.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 266.546 934.59 267.694 ;
      VIA 933.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 256.466 934.59 257.614 ;
      VIA 933.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 933.556 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.556 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.428 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.3 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.172 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 933.044 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  932.45 14.546 934.59 15.694 ;
      VIA 933.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 933.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 609.266 889.79 610.414 ;
      VIA 888.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 599.186 889.79 600.334 ;
      VIA 888.976 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 589.106 889.79 590.254 ;
      VIA 888.976 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 347.186 889.79 348.334 ;
      VIA 888.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 337.106 889.79 338.254 ;
      VIA 888.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 327.026 889.79 328.174 ;
      VIA 888.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 316.946 889.79 318.094 ;
      VIA 888.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 306.866 889.79 308.014 ;
      VIA 888.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 296.786 889.79 297.934 ;
      VIA 888.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 286.706 889.79 287.854 ;
      VIA 888.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 276.626 889.79 277.774 ;
      VIA 888.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 266.546 889.79 267.694 ;
      VIA 888.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 256.466 889.79 257.614 ;
      VIA 888.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 888.556 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.556 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.428 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.3 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.172 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 888.044 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  887.65 14.546 889.79 15.694 ;
      VIA 888.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 888.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 609.266 844.99 610.414 ;
      VIA 844.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 599.186 844.99 600.334 ;
      VIA 844.176 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 589.106 844.99 590.254 ;
      VIA 844.176 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 347.186 844.99 348.334 ;
      VIA 844.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 337.106 844.99 338.254 ;
      VIA 844.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 327.026 844.99 328.174 ;
      VIA 844.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 316.946 844.99 318.094 ;
      VIA 844.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 306.866 844.99 308.014 ;
      VIA 844.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 296.786 844.99 297.934 ;
      VIA 844.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 286.706 844.99 287.854 ;
      VIA 844.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 276.626 844.99 277.774 ;
      VIA 844.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 266.546 844.99 267.694 ;
      VIA 844.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 256.466 844.99 257.614 ;
      VIA 844.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 844.456 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.456 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.328 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.2 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 844.072 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 843.944 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  842.85 14.546 844.99 15.694 ;
      VIA 844.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 844.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 843.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 609.266 800.19 610.414 ;
      VIA 799.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 599.186 800.19 600.334 ;
      VIA 799.376 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 589.106 800.19 590.254 ;
      VIA 799.376 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 347.186 800.19 348.334 ;
      VIA 799.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 337.106 800.19 338.254 ;
      VIA 799.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 327.026 800.19 328.174 ;
      VIA 799.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 316.946 800.19 318.094 ;
      VIA 799.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 306.866 800.19 308.014 ;
      VIA 799.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 296.786 800.19 297.934 ;
      VIA 799.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 286.706 800.19 287.854 ;
      VIA 799.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 276.626 800.19 277.774 ;
      VIA 799.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 266.546 800.19 267.694 ;
      VIA 799.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 256.466 800.19 257.614 ;
      VIA 799.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 799.456 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.456 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.328 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.2 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 799.072 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 798.944 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  798.05 14.546 800.19 15.694 ;
      VIA 799.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 798.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 799.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 609.266 755.39 610.414 ;
      VIA 754.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 599.186 755.39 600.334 ;
      VIA 754.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 589.106 755.39 590.254 ;
      VIA 754.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 347.186 755.39 348.334 ;
      VIA 754.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 337.106 755.39 338.254 ;
      VIA 754.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 327.026 755.39 328.174 ;
      VIA 754.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 316.946 755.39 318.094 ;
      VIA 754.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 306.866 755.39 308.014 ;
      VIA 754.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 296.786 755.39 297.934 ;
      VIA 754.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 286.706 755.39 287.854 ;
      VIA 754.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 276.626 755.39 277.774 ;
      VIA 754.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 266.546 755.39 267.694 ;
      VIA 754.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 256.466 755.39 257.614 ;
      VIA 754.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 754.456 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.456 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.328 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.2 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 754.072 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 753.944 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  753.25 14.546 755.39 15.694 ;
      VIA 754.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 754.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 609.266 710.59 610.414 ;
      VIA 709.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 599.186 710.59 600.334 ;
      VIA 709.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 589.106 710.59 590.254 ;
      VIA 709.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 347.186 710.59 348.334 ;
      VIA 709.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 337.106 710.59 338.254 ;
      VIA 709.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 327.026 710.59 328.174 ;
      VIA 709.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 316.946 710.59 318.094 ;
      VIA 709.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 306.866 710.59 308.014 ;
      VIA 709.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 296.786 710.59 297.934 ;
      VIA 709.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 286.706 710.59 287.854 ;
      VIA 709.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 276.626 710.59 277.774 ;
      VIA 709.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 266.546 710.59 267.694 ;
      VIA 709.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 256.466 710.59 257.614 ;
      VIA 709.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 709.456 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.456 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.328 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.2 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 709.072 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 708.944 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  708.45 14.546 710.59 15.694 ;
      VIA 709.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 709.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 609.266 665.79 610.414 ;
      VIA 664.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 599.186 665.79 600.334 ;
      VIA 664.976 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 589.106 665.79 590.254 ;
      VIA 664.976 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 347.186 665.79 348.334 ;
      VIA 664.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 337.106 665.79 338.254 ;
      VIA 664.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 327.026 665.79 328.174 ;
      VIA 664.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 316.946 665.79 318.094 ;
      VIA 664.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 306.866 665.79 308.014 ;
      VIA 664.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 296.786 665.79 297.934 ;
      VIA 664.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 286.706 665.79 287.854 ;
      VIA 664.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 276.626 665.79 277.774 ;
      VIA 664.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 266.546 665.79 267.694 ;
      VIA 664.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 256.466 665.79 257.614 ;
      VIA 664.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 665.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 665.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 664.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  663.65 14.546 665.79 15.694 ;
      VIA 664.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 664.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 609.266 620.99 610.414 ;
      VIA 620.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 599.186 620.99 600.334 ;
      VIA 620.176 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 589.106 620.99 590.254 ;
      VIA 620.176 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 347.186 620.99 348.334 ;
      VIA 620.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 337.106 620.99 338.254 ;
      VIA 620.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 327.026 620.99 328.174 ;
      VIA 620.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 316.946 620.99 318.094 ;
      VIA 620.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 306.866 620.99 308.014 ;
      VIA 620.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 296.786 620.99 297.934 ;
      VIA 620.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 286.706 620.99 287.854 ;
      VIA 620.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 276.626 620.99 277.774 ;
      VIA 620.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 266.546 620.99 267.694 ;
      VIA 620.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 256.466 620.99 257.614 ;
      VIA 620.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 620.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 620.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 619.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  618.85 14.546 620.99 15.694 ;
      VIA 620.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 620.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 619.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 609.266 576.19 610.414 ;
      VIA 575.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 599.186 576.19 600.334 ;
      VIA 575.376 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 589.106 576.19 590.254 ;
      VIA 575.376 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 347.186 576.19 348.334 ;
      VIA 575.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 337.106 576.19 338.254 ;
      VIA 575.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 327.026 576.19 328.174 ;
      VIA 575.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 316.946 576.19 318.094 ;
      VIA 575.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 306.866 576.19 308.014 ;
      VIA 575.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 296.786 576.19 297.934 ;
      VIA 575.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 286.706 576.19 287.854 ;
      VIA 575.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 276.626 576.19 277.774 ;
      VIA 575.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 266.546 576.19 267.694 ;
      VIA 575.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 256.466 576.19 257.614 ;
      VIA 575.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 14.546 576.19 15.694 ;
      VIA 575.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 609.266 531.39 610.414 ;
      VIA 530.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 599.186 531.39 600.334 ;
      VIA 530.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 589.106 531.39 590.254 ;
      VIA 530.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 579.026 531.39 580.174 ;
      VIA 530.576 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 568.946 531.39 570.094 ;
      VIA 530.576 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 558.866 531.39 560.014 ;
      VIA 530.576 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 548.786 531.39 549.934 ;
      VIA 530.576 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 538.706 531.39 539.854 ;
      VIA 530.576 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 528.626 531.39 529.774 ;
      VIA 530.576 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 518.546 531.39 519.694 ;
      VIA 530.576 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 508.466 531.39 509.614 ;
      VIA 530.576 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 498.386 531.39 499.534 ;
      VIA 530.576 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 488.306 531.39 489.454 ;
      VIA 530.576 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 478.226 531.39 479.374 ;
      VIA 530.576 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 468.146 531.39 469.294 ;
      VIA 530.576 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 458.066 531.39 459.214 ;
      VIA 530.576 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 447.986 531.39 449.134 ;
      VIA 530.576 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 437.906 531.39 439.054 ;
      VIA 530.576 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 427.826 531.39 428.974 ;
      VIA 530.576 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 417.746 531.39 418.894 ;
      VIA 530.576 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 407.666 531.39 408.814 ;
      VIA 530.576 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 397.586 531.39 398.734 ;
      VIA 530.576 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 387.506 531.39 388.654 ;
      VIA 530.576 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 377.426 531.39 378.574 ;
      VIA 530.576 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 367.346 531.39 368.494 ;
      VIA 530.576 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 357.266 531.39 358.414 ;
      VIA 530.576 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 347.186 531.39 348.334 ;
      VIA 530.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 337.106 531.39 338.254 ;
      VIA 530.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 327.026 531.39 328.174 ;
      VIA 530.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 316.946 531.39 318.094 ;
      VIA 530.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 306.866 531.39 308.014 ;
      VIA 530.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 296.786 531.39 297.934 ;
      VIA 530.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 286.706 531.39 287.854 ;
      VIA 530.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 276.626 531.39 277.774 ;
      VIA 530.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 266.546 531.39 267.694 ;
      VIA 530.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 256.466 531.39 257.614 ;
      VIA 530.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 246.386 531.39 247.534 ;
      VIA 530.576 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 236.306 531.39 237.454 ;
      VIA 530.576 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 226.226 531.39 227.374 ;
      VIA 530.576 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 216.146 531.39 217.294 ;
      VIA 530.576 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 206.066 531.39 207.214 ;
      VIA 530.576 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 195.986 531.39 197.134 ;
      VIA 530.576 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 185.906 531.39 187.054 ;
      VIA 530.576 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 175.826 531.39 176.974 ;
      VIA 530.576 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 165.746 531.39 166.894 ;
      VIA 530.576 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 155.666 531.39 156.814 ;
      VIA 530.576 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 145.586 531.39 146.734 ;
      VIA 530.576 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 135.506 531.39 136.654 ;
      VIA 530.576 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 125.426 531.39 126.574 ;
      VIA 530.576 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 115.346 531.39 116.494 ;
      VIA 530.576 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 105.266 531.39 106.414 ;
      VIA 530.576 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 95.186 531.39 96.334 ;
      VIA 530.576 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 85.106 531.39 86.254 ;
      VIA 530.576 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 75.026 531.39 76.174 ;
      VIA 530.576 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 64.946 531.39 66.094 ;
      VIA 530.576 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 54.866 531.39 56.014 ;
      VIA 530.576 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 44.786 531.39 45.934 ;
      VIA 530.576 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 34.706 531.39 35.854 ;
      VIA 530.576 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 24.626 531.39 25.774 ;
      VIA 530.576 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 14.546 531.39 15.694 ;
      VIA 530.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 609.266 486.59 610.414 ;
      VIA 485.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 599.186 486.59 600.334 ;
      VIA 485.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 589.106 486.59 590.254 ;
      VIA 485.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 579.026 486.59 580.174 ;
      VIA 485.776 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 568.946 486.59 570.094 ;
      VIA 485.776 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 558.866 486.59 560.014 ;
      VIA 485.776 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 548.786 486.59 549.934 ;
      VIA 485.776 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 538.706 486.59 539.854 ;
      VIA 485.776 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 528.626 486.59 529.774 ;
      VIA 485.776 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 518.546 486.59 519.694 ;
      VIA 485.776 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 508.466 486.59 509.614 ;
      VIA 485.776 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 498.386 486.59 499.534 ;
      VIA 485.776 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 488.306 486.59 489.454 ;
      VIA 485.776 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 478.226 486.59 479.374 ;
      VIA 485.776 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 468.146 486.59 469.294 ;
      VIA 485.776 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 458.066 486.59 459.214 ;
      VIA 485.776 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 447.986 486.59 449.134 ;
      VIA 485.776 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 437.906 486.59 439.054 ;
      VIA 485.776 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 427.826 486.59 428.974 ;
      VIA 485.776 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 417.746 486.59 418.894 ;
      VIA 485.776 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 407.666 486.59 408.814 ;
      VIA 485.776 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 397.586 486.59 398.734 ;
      VIA 485.776 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 387.506 486.59 388.654 ;
      VIA 485.776 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 377.426 486.59 378.574 ;
      VIA 485.776 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 367.346 486.59 368.494 ;
      VIA 485.776 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 357.266 486.59 358.414 ;
      VIA 485.776 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 347.186 486.59 348.334 ;
      VIA 485.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 337.106 486.59 338.254 ;
      VIA 485.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 327.026 486.59 328.174 ;
      VIA 485.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 316.946 486.59 318.094 ;
      VIA 485.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 306.866 486.59 308.014 ;
      VIA 485.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 296.786 486.59 297.934 ;
      VIA 485.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 286.706 486.59 287.854 ;
      VIA 485.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 276.626 486.59 277.774 ;
      VIA 485.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 266.546 486.59 267.694 ;
      VIA 485.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 256.466 486.59 257.614 ;
      VIA 485.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 246.386 486.59 247.534 ;
      VIA 485.776 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 236.306 486.59 237.454 ;
      VIA 485.776 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 226.226 486.59 227.374 ;
      VIA 485.776 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 216.146 486.59 217.294 ;
      VIA 485.776 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 206.066 486.59 207.214 ;
      VIA 485.776 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 195.986 486.59 197.134 ;
      VIA 485.776 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 185.906 486.59 187.054 ;
      VIA 485.776 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 175.826 486.59 176.974 ;
      VIA 485.776 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 165.746 486.59 166.894 ;
      VIA 485.776 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 155.666 486.59 156.814 ;
      VIA 485.776 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 145.586 486.59 146.734 ;
      VIA 485.776 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 135.506 486.59 136.654 ;
      VIA 485.776 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 125.426 486.59 126.574 ;
      VIA 485.776 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 115.346 486.59 116.494 ;
      VIA 485.776 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 105.266 486.59 106.414 ;
      VIA 485.776 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 95.186 486.59 96.334 ;
      VIA 485.776 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 85.106 486.59 86.254 ;
      VIA 485.776 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 75.026 486.59 76.174 ;
      VIA 485.776 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 64.946 486.59 66.094 ;
      VIA 485.776 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 54.866 486.59 56.014 ;
      VIA 485.776 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 44.786 486.59 45.934 ;
      VIA 485.776 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 34.706 486.59 35.854 ;
      VIA 485.776 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 24.626 486.59 25.774 ;
      VIA 485.776 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 14.546 486.59 15.694 ;
      VIA 485.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 609.266 441.79 610.414 ;
      VIA 440.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 599.186 441.79 600.334 ;
      VIA 440.976 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 589.106 441.79 590.254 ;
      VIA 440.976 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 347.186 441.79 348.334 ;
      VIA 440.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 337.106 441.79 338.254 ;
      VIA 440.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 327.026 441.79 328.174 ;
      VIA 440.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 316.946 441.79 318.094 ;
      VIA 440.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 306.866 441.79 308.014 ;
      VIA 440.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 296.786 441.79 297.934 ;
      VIA 440.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 286.706 441.79 287.854 ;
      VIA 440.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 276.626 441.79 277.774 ;
      VIA 440.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 266.546 441.79 267.694 ;
      VIA 440.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 256.466 441.79 257.614 ;
      VIA 440.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 14.546 441.79 15.694 ;
      VIA 440.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 609.266 396.99 610.414 ;
      VIA 396.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 599.186 396.99 600.334 ;
      VIA 396.176 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 589.106 396.99 590.254 ;
      VIA 396.176 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 347.186 396.99 348.334 ;
      VIA 396.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 337.106 396.99 338.254 ;
      VIA 396.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 327.026 396.99 328.174 ;
      VIA 396.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 316.946 396.99 318.094 ;
      VIA 396.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 306.866 396.99 308.014 ;
      VIA 396.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 296.786 396.99 297.934 ;
      VIA 396.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 286.706 396.99 287.854 ;
      VIA 396.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 276.626 396.99 277.774 ;
      VIA 396.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 266.546 396.99 267.694 ;
      VIA 396.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 256.466 396.99 257.614 ;
      VIA 396.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 14.546 396.99 15.694 ;
      VIA 396.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 609.266 352.19 610.414 ;
      VIA 351.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 599.186 352.19 600.334 ;
      VIA 351.376 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 589.106 352.19 590.254 ;
      VIA 351.376 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 347.186 352.19 348.334 ;
      VIA 351.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 337.106 352.19 338.254 ;
      VIA 351.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 327.026 352.19 328.174 ;
      VIA 351.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 316.946 352.19 318.094 ;
      VIA 351.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 306.866 352.19 308.014 ;
      VIA 351.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 296.786 352.19 297.934 ;
      VIA 351.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 286.706 352.19 287.854 ;
      VIA 351.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 276.626 352.19 277.774 ;
      VIA 351.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 266.546 352.19 267.694 ;
      VIA 351.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 256.466 352.19 257.614 ;
      VIA 351.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 14.546 352.19 15.694 ;
      VIA 351.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 609.266 307.39 610.414 ;
      VIA 306.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 599.186 307.39 600.334 ;
      VIA 306.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 589.106 307.39 590.254 ;
      VIA 306.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 347.186 307.39 348.334 ;
      VIA 306.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 337.106 307.39 338.254 ;
      VIA 306.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 327.026 307.39 328.174 ;
      VIA 306.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 316.946 307.39 318.094 ;
      VIA 306.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 306.866 307.39 308.014 ;
      VIA 306.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 296.786 307.39 297.934 ;
      VIA 306.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 286.706 307.39 287.854 ;
      VIA 306.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 276.626 307.39 277.774 ;
      VIA 306.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 266.546 307.39 267.694 ;
      VIA 306.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 256.466 307.39 257.614 ;
      VIA 306.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 14.546 307.39 15.694 ;
      VIA 306.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 609.266 262.59 610.414 ;
      VIA 261.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 599.186 262.59 600.334 ;
      VIA 261.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 589.106 262.59 590.254 ;
      VIA 261.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 347.186 262.59 348.334 ;
      VIA 261.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 337.106 262.59 338.254 ;
      VIA 261.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 327.026 262.59 328.174 ;
      VIA 261.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 316.946 262.59 318.094 ;
      VIA 261.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 306.866 262.59 308.014 ;
      VIA 261.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 296.786 262.59 297.934 ;
      VIA 261.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 286.706 262.59 287.854 ;
      VIA 261.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 276.626 262.59 277.774 ;
      VIA 261.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 266.546 262.59 267.694 ;
      VIA 261.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 256.466 262.59 257.614 ;
      VIA 261.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 14.546 262.59 15.694 ;
      VIA 261.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 609.266 217.79 610.414 ;
      VIA 216.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 599.186 217.79 600.334 ;
      VIA 216.976 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 589.106 217.79 590.254 ;
      VIA 216.976 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 347.186 217.79 348.334 ;
      VIA 216.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 337.106 217.79 338.254 ;
      VIA 216.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 327.026 217.79 328.174 ;
      VIA 216.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 316.946 217.79 318.094 ;
      VIA 216.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 306.866 217.79 308.014 ;
      VIA 216.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 296.786 217.79 297.934 ;
      VIA 216.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 286.706 217.79 287.854 ;
      VIA 216.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 276.626 217.79 277.774 ;
      VIA 216.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 266.546 217.79 267.694 ;
      VIA 216.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 256.466 217.79 257.614 ;
      VIA 216.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 14.546 217.79 15.694 ;
      VIA 216.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 609.266 172.99 610.414 ;
      VIA 172.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 599.186 172.99 600.334 ;
      VIA 172.176 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 589.106 172.99 590.254 ;
      VIA 172.176 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 347.186 172.99 348.334 ;
      VIA 172.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 337.106 172.99 338.254 ;
      VIA 172.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 327.026 172.99 328.174 ;
      VIA 172.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 316.946 172.99 318.094 ;
      VIA 172.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 306.866 172.99 308.014 ;
      VIA 172.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 296.786 172.99 297.934 ;
      VIA 172.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 286.706 172.99 287.854 ;
      VIA 172.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 276.626 172.99 277.774 ;
      VIA 172.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 266.546 172.99 267.694 ;
      VIA 172.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 256.466 172.99 257.614 ;
      VIA 172.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 14.546 172.99 15.694 ;
      VIA 172.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 609.266 128.19 610.414 ;
      VIA 127.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 599.186 128.19 600.334 ;
      VIA 127.376 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 589.106 128.19 590.254 ;
      VIA 127.376 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 347.186 128.19 348.334 ;
      VIA 127.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 337.106 128.19 338.254 ;
      VIA 127.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 327.026 128.19 328.174 ;
      VIA 127.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 316.946 128.19 318.094 ;
      VIA 127.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 306.866 128.19 308.014 ;
      VIA 127.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 296.786 128.19 297.934 ;
      VIA 127.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 286.706 128.19 287.854 ;
      VIA 127.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 276.626 128.19 277.774 ;
      VIA 127.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 266.546 128.19 267.694 ;
      VIA 127.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 256.466 128.19 257.614 ;
      VIA 127.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 14.546 128.19 15.694 ;
      VIA 127.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 609.266 83.39 610.414 ;
      VIA 82.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 599.186 83.39 600.334 ;
      VIA 82.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 589.106 83.39 590.254 ;
      VIA 82.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 347.186 83.39 348.334 ;
      VIA 82.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 337.106 83.39 338.254 ;
      VIA 82.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 327.026 83.39 328.174 ;
      VIA 82.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 316.946 83.39 318.094 ;
      VIA 82.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 306.866 83.39 308.014 ;
      VIA 82.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 296.786 83.39 297.934 ;
      VIA 82.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 286.706 83.39 287.854 ;
      VIA 82.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 276.626 83.39 277.774 ;
      VIA 82.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 266.546 83.39 267.694 ;
      VIA 82.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 256.466 83.39 257.614 ;
      VIA 82.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 14.546 83.39 15.694 ;
      VIA 82.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 609.266 38.59 610.414 ;
      VIA 37.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 599.186 38.59 600.334 ;
      VIA 37.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 589.106 38.59 590.254 ;
      VIA 37.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 347.186 38.59 348.334 ;
      VIA 37.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 337.106 38.59 338.254 ;
      VIA 37.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 327.026 38.59 328.174 ;
      VIA 37.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 316.946 38.59 318.094 ;
      VIA 37.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 306.866 38.59 308.014 ;
      VIA 37.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 296.786 38.59 297.934 ;
      VIA 37.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 286.706 38.59 287.854 ;
      VIA 37.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 276.626 38.59 277.774 ;
      VIA 37.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 266.546 38.59 267.694 ;
      VIA 37.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 256.466 38.59 257.614 ;
      VIA 37.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 14.546 38.59 15.694 ;
      VIA 37.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 12.856 590.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 590.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 590.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 590.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 590.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 589.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 589.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 589.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 589.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 589.296 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 589.106 13.39 590.254 ;
      VIA 12.576 590.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 590.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 590.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 590.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 590.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 589.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 589.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 589.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 589.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 589.68 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 579.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 579.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 579.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 579.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 579.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 579.216 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 579.026 13.39 580.174 ;
      VIA 12.576 579.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 579.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 579.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 579.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 579.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 579.6 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 569.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 569.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 569.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 569.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 569.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 569.136 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 568.946 13.39 570.094 ;
      VIA 12.576 569.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 569.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 569.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 569.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 569.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 569.52 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 559.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 559.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 559.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 559.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 559.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 559.056 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 558.866 13.39 560.014 ;
      VIA 12.576 559.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 559.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 559.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 559.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 559.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 559.44 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 549.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 549.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 549.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 549.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 549.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 549.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 549.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 549.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 549.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 549.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 548.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 548.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 548.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 548.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 548.976 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 548.786 13.39 549.934 ;
      VIA 12.576 549.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 549.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 549.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 549.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 549.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 549.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 549.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 549.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 549.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 548.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 548.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 548.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 548.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 548.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 549.36 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 539.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 539.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 539.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 539.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 539.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 539.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 539.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 539.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 539.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 539.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 538.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 538.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 538.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 538.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 538.896 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 538.706 13.39 539.854 ;
      VIA 12.576 539.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 539.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 539.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 539.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 539.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 539.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 539.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 539.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 539.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 538.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 538.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 538.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 538.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 538.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 539.28 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 529.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 529.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 529.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 529.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 529.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 529.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 529.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 529.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 529.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 529.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 529.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 529.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 529.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 529.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 529.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 529.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 529.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 529.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 529.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 529.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 529.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 529.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 529.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 529.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 529.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 528.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 528.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 528.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 528.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 528.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 528.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 528.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 528.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 528.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 528.816 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 528.626 13.39 529.774 ;
      VIA 12.576 529.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 529.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 529.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 529.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 529.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 529.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 529.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 529.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 529.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 529.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 529.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 529.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 529.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 529.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 529.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 529.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 529.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 529.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 529.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 529.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 528.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 528.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 528.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 528.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 528.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 528.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 528.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 528.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 528.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 528.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 529.2 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 519.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 519.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 519.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 519.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 519.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 519.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 519.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 519.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 519.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 519.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 519.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 519.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 519.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 519.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 519.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 519.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 519.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 519.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 519.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 519.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 518.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 518.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 518.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 518.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 518.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 518.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 518.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 518.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 518.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 518.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 518.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 518.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 518.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 518.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 518.736 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 518.546 13.39 519.694 ;
      VIA 12.576 519.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 519.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 519.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 519.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 519.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 519.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 519.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 519.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 519.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 519.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 519.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 519.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 519.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 519.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 519.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 519.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 519.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 519.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 519.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 519.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 518.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 518.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 518.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 518.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 518.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 518.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 518.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 518.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 518.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 518.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 518.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 518.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 518.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 518.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 518.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 519.12 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 509.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 509.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 509.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 509.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 509.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 509.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 509.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 509.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 509.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 509.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 509.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 509.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 509.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 509.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 509.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 509.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 509.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 509.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 509.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 509.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 508.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 508.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 508.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 508.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 508.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 508.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 508.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 508.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 508.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 508.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 508.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 508.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 508.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 508.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 508.656 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 508.466 13.39 509.614 ;
      VIA 12.576 509.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 509.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 509.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 509.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 509.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 509.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 509.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 509.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 509.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 509.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 509.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 509.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 509.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 509.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 509.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 509.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 509.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 509.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 509.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 509.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 508.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 508.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 508.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 508.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 508.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 508.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 508.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 508.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 508.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 508.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 508.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 508.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 508.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 508.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 508.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 509.04 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 499.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 499.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 499.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 499.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 499.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 499.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 499.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 499.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 499.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 499.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 499.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 499.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 499.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 499.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 499.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 498.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 498.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 498.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 498.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 498.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 498.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 498.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 498.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 498.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 498.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 498.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 498.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 498.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 498.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 498.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 498.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 498.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 498.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 498.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 498.576 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 498.386 13.39 499.534 ;
      VIA 12.576 499.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 499.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 499.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 499.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 499.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 499.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 499.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 499.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 499.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 499.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 499.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 499.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 499.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 499.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 499.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 498.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 498.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 498.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 498.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 498.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 498.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 498.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 498.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 498.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 498.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 498.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 498.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 498.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 498.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 498.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 498.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 498.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 498.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 498.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 498.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 498.96 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 489.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 489.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 489.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 489.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 489.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 489.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 489.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 489.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 489.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 489.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 489.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 489.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 489.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 489.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 489.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 488.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 488.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 488.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 488.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 488.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 488.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 488.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 488.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 488.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 488.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 488.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 488.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 488.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 488.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 488.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 488.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 488.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 488.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 488.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 488.496 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 488.306 13.39 489.454 ;
      VIA 12.576 489.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 489.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 489.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 489.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 489.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 489.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 489.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 489.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 489.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 489.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 489.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 489.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 489.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 489.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 489.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 488.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 488.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 488.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 488.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 488.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 488.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 488.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 488.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 488.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 488.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 488.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 488.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 488.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 488.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 488.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 488.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 488.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 488.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 488.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 488.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 488.88 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 479.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 479.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 479.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 479.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 479.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 479.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 479.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 479.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 479.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 479.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 478.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 478.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 478.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 478.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 478.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 478.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 478.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 478.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 478.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 478.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 478.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 478.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 478.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 478.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 478.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 478.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 478.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 478.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 478.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 478.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 478.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 478.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 478.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 478.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 478.416 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 478.226 13.39 479.374 ;
      VIA 12.576 479.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 479.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 479.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 479.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 479.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 479.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 479.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 479.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 479.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 479.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 478.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 478.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 478.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 478.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 478.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 478.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 478.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 478.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 478.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 478.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 478.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 478.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 478.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 478.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 478.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 478.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 478.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 478.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 478.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 478.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 478.8 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 469.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 469.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 469.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 469.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 469.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 468.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 468.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 468.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 468.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 468.336 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 468.146 13.39 469.294 ;
      VIA 12.576 469.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 469.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 469.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 469.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 469.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 468.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 468.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 468.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 468.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 468.72 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 459.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 459.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 459.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 459.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 459.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 458.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 458.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 458.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 458.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 458.256 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 458.066 13.39 459.214 ;
      VIA 12.576 459.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 459.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 459.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 459.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 459.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 458.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 458.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 458.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 458.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 458.64 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 448.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 448.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 448.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 448.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 448.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 448.176 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 447.986 13.39 449.134 ;
      VIA 12.576 448.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 448.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 448.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 448.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 448.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 448.56 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 438.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 438.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 438.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 438.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 438.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 438.096 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 437.906 13.39 439.054 ;
      VIA 12.576 438.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 438.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 438.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 438.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 438.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 438.48 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 428.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 428.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 428.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 428.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 428.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 428.016 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 427.826 13.39 428.974 ;
      VIA 12.576 428.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 428.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 428.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 428.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 428.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 428.4 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 418.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 418.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 418.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 418.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 418.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 418.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 418.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 418.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 418.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 418.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 417.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 417.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 417.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 417.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 417.936 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 417.746 13.39 418.894 ;
      VIA 12.576 418.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 418.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 418.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 418.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 418.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 418.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 418.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 418.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 418.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 417.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 417.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 417.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 417.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 417.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 418.32 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 408.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 408.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 408.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 408.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 408.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 408.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 408.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 408.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 408.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 408.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 408.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 408.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 408.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 408.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 408.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 408.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 408.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 408.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 408.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 408.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 408.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 408.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 408.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 408.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 408.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 407.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 407.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 407.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 407.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 407.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 407.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 407.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 407.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 407.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 407.856 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 407.666 13.39 408.814 ;
      VIA 12.576 408.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 408.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 408.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 408.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 408.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 408.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 408.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 408.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 408.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 408.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 408.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 408.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 408.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 408.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 408.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 408.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 408.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 408.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 408.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 408.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 407.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 407.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 407.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 407.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 407.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 407.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 407.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 407.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 407.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 407.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 408.24 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 398.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 398.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 398.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 398.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 398.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 398.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 398.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 398.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 398.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 398.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 398.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 398.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 398.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 398.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 398.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 398.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 398.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 398.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 398.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 398.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 398.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 398.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 398.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 398.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 398.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 397.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 397.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 397.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 397.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 397.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 397.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 397.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 397.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 397.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 397.776 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 397.586 13.39 398.734 ;
      VIA 12.576 398.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 398.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 398.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 398.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 398.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 398.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 398.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 398.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 398.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 398.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 398.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 398.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 398.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 398.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 398.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 398.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 398.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 398.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 398.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 398.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 397.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 397.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 397.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 397.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 397.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 397.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 397.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 397.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 397.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 397.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 398.16 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 388.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 388.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 388.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 388.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 388.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 388.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 388.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 388.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 388.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 388.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 388.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 388.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 388.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 388.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 388.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 388.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 388.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 388.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 388.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 388.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 387.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 387.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 387.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 387.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 387.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 387.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 387.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 387.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 387.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 387.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 387.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 387.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 387.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 387.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 387.696 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 387.506 13.39 388.654 ;
      VIA 12.576 388.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 388.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 388.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 388.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 388.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 388.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 388.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 388.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 388.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 388.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 388.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 388.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 388.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 388.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 388.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 388.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 388.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 388.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 388.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 388.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 387.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 387.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 387.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 387.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 387.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 387.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 387.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 387.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 387.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 387.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 387.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 387.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 387.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 387.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 387.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 388.08 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 378.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 378.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 378.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 378.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 378.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 378.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 378.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 378.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 378.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 378.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 378.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 378.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 378.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 378.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 378.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 378 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 378 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 378 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 378 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 378 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 377.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 377.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 377.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 377.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 377.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 377.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 377.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 377.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 377.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 377.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 377.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 377.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 377.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 377.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 377.616 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 377.426 13.39 378.574 ;
      VIA 12.576 378.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 378.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 378.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 378.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 378.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 378.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 378.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 378.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 378.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 378.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 378.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 378.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 378.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 378.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 378.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 378 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 378 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 378 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 378 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 378 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 377.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 377.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 377.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 377.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 377.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 377.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 377.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 377.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 377.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 377.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 377.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 377.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 377.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 377.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 377.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 378 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 368.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 368.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 368.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 368.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 368.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 368.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 368.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 368.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 368.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 368.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 368.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 368.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 368.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 368.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 368.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 367.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 367.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 367.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 367.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 367.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 367.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 367.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 367.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 367.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 367.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 367.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 367.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 367.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 367.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 367.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 367.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 367.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 367.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 367.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 367.536 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 367.346 13.39 368.494 ;
      VIA 12.576 368.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 368.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 368.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 368.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 368.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 368.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 368.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 368.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 368.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 368.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 368.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 368.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 368.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 368.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 368.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 367.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 367.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 367.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 367.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 367.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 367.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 367.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 367.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 367.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 367.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 367.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 367.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 367.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 367.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 367.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 367.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 367.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 367.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 367.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 367.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 367.92 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 358.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 358.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 358.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 358.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 358.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 358.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 358.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 358.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 358.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 358.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 357.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 357.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 357.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 357.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 357.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 357.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 357.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 357.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 357.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 357.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 357.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 357.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 357.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 357.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 357.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 357.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 357.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 357.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 357.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 357.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 357.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 357.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 357.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 357.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 357.456 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 357.266 13.39 358.414 ;
      VIA 12.576 358.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 358.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 358.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 358.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 358.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 358.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 358.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 358.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 358.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 358.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 357.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 357.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 357.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 357.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 357.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 357.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 357.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 357.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 357.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 357.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 357.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 357.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 357.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 357.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 357.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 357.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 357.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 357.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 357.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 357.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 357.84 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 348.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 348.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 348.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 348.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 348.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 348.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 348.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 348.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 348.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 348.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 347.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 347.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 347.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 347.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 347.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 347.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 347.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 347.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 347.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 347.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 347.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 347.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 347.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 347.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 347.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 347.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 347.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 347.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 347.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 347.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 347.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 347.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 347.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 347.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 347.376 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 347.186 13.39 348.334 ;
      VIA 12.576 348.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 348.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 348.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 348.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 348.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 348.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 348.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 348.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 348.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 348.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 347.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 347.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 347.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 347.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 347.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 347.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 347.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 347.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 347.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 347.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 347.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 347.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 347.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 347.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 347.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 347.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 347.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 347.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 347.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 347.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 347.76 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 257.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 257.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 257.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 257.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 257.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 257.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 257.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 257.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 257.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 257.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 257.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 257.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 257.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 257.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 257.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 257.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 257.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 257.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 257.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 257.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 256.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 256.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 256.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 256.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 256.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 256.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 256.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 256.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 256.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 256.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 256.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 256.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 256.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 256.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 256.656 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 256.466 13.39 257.614 ;
      VIA 12.576 257.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 257.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 257.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 257.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 257.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 257.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 257.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 257.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 257.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 257.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 257.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 257.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 257.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 257.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 257.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 257.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 257.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 257.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 257.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 257.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 256.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 256.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 256.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 256.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 256.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 256.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 256.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 256.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 256.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 256.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 256.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 256.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 256.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 256.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 256.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 257.04 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 247.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 247.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 247.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 247.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 247.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 247.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 247.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 247.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 247.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 247.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 247.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 247.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 247.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 247.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 247.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 246.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 246.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 246.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 246.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 246.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 246.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 246.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 246.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 246.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 246.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 246.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 246.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 246.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 246.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 246.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 246.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 246.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 246.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 246.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 246.576 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 246.386 13.39 247.534 ;
      VIA 12.576 247.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 247.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 247.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 247.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 247.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 247.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 247.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 247.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 247.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 247.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 247.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 247.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 247.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 247.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 247.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 246.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 246.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 246.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 246.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 246.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 246.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 246.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 246.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 246.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 246.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 246.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 246.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 246.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 246.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 246.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 246.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 246.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 246.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 246.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 246.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 246.96 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 237.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 237.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 237.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 237.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 237.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 237.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 237.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 237.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 237.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 237.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 237.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 237.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 237.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 237.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 237.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 236.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 236.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 236.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 236.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 236.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 236.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 236.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 236.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 236.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 236.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 236.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 236.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 236.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 236.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 236.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 236.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 236.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 236.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 236.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 236.496 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 236.306 13.39 237.454 ;
      VIA 12.576 237.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 237.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 237.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 237.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 237.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 237.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 237.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 237.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 237.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 237.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 237.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 237.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 237.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 237.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 237.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 236.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 236.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 236.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 236.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 236.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 236.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 236.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 236.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 236.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 236.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 236.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 236.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 236.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 236.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 236.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 236.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 236.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 236.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 236.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 236.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 236.88 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 227.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 227.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 227.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 227.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 227.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 227.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 227.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 227.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 227.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 227.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 226.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 226.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 226.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 226.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 226.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 226.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 226.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 226.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 226.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 226.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 226.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 226.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 226.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 226.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 226.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 226.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 226.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 226.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 226.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 226.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 226.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 226.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 226.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 226.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 226.416 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 226.226 13.39 227.374 ;
      VIA 12.576 227.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 227.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 227.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 227.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 227.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 227.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 227.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 227.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 227.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 227.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 226.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 226.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 226.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 226.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 226.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 226.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 226.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 226.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 226.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 226.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 226.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 226.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 226.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 226.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 226.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 226.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 226.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 226.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 226.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 226.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 226.8 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 217.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 217.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 217.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 217.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 217.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 216.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 216.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 216.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 216.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 216.336 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 216.146 13.39 217.294 ;
      VIA 12.576 217.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 217.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 217.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 217.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 217.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 216.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 216.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 216.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 216.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 216.72 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 207.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 207.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 207.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 207.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 207.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 206.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 206.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 206.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 206.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 206.256 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 206.066 13.39 207.214 ;
      VIA 12.576 207.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 207.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 207.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 207.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 207.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 206.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 206.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 206.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 206.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 206.64 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 196.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 196.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 196.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 196.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 196.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 196.176 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 195.986 13.39 197.134 ;
      VIA 12.576 196.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 196.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 196.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 196.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 196.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 196.56 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 186.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 186.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 186.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 186.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 186.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 186.096 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 185.906 13.39 187.054 ;
      VIA 12.576 186.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 186.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 186.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 186.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 186.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 186.48 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 176.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 176.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 176.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 176.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 176.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 176.016 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 175.826 13.39 176.974 ;
      VIA 12.576 176.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 176.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 176.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 176.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 176.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 176.4 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 166.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 166.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 166.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 166.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 166.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 166.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 166.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 166.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 166.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 166.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 165.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 165.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 165.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 165.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 165.936 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 165.746 13.39 166.894 ;
      VIA 12.576 166.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 166.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 166.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 166.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 166.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 166.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 166.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 166.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 166.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 165.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 165.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 165.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 165.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 165.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 166.32 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 156.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 156.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 156.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 156.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 156.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 156.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 156.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 156.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 156.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 156.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 156.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 156.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 156.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 156.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 156.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 156.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 156.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 156.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 156.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 156.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 156.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 156.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 156.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 156.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 156.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 155.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 155.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 155.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 155.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 155.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 155.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 155.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 155.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 155.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 155.856 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 155.666 13.39 156.814 ;
      VIA 12.576 156.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 156.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 156.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 156.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 156.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 156.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 156.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 156.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 156.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 156.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 156.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 156.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 156.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 156.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 156.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 156.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 156.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 156.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 156.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 156.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 155.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 155.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 155.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 155.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 155.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 155.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 155.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 155.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 155.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 155.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 156.24 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 146.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 146.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 146.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 146.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 146.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 146.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 146.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 146.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 146.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 146.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 146.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 146.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 146.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 146.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 146.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 146.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 146.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 146.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 146.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 146.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 146.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 146.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 146.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 146.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 146.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 145.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 145.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 145.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 145.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 145.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 145.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 145.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 145.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 145.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 145.776 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 145.586 13.39 146.734 ;
      VIA 12.576 146.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 146.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 146.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 146.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 146.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 146.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 146.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 146.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 146.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 146.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 146.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 146.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 146.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 146.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 146.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 146.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 146.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 146.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 146.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 146.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 145.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 145.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 145.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 145.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 145.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 145.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 145.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 145.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 145.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 145.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 146.16 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 136.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 136.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 136.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 136.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 136.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 136.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 136.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 136.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 136.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 136.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 136.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 136.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 136.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 136.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 136.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 136.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 136.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 136.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 136.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 136.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 135.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 135.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 135.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 135.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 135.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 135.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 135.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 135.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 135.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 135.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 135.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 135.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 135.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 135.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 135.696 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 135.506 13.39 136.654 ;
      VIA 12.576 136.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 136.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 136.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 136.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 136.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 136.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 136.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 136.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 136.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 136.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 136.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 136.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 136.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 136.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 136.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 136.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 136.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 136.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 136.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 136.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 135.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 135.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 135.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 135.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 135.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 135.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 135.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 135.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 135.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 135.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 135.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 135.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 135.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 135.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 135.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 136.08 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 126.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 126.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 126.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 126.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 126.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 126.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 126.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 126.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 126.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 126.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 126.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 126.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 126.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 126.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 126.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 126 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 126 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 126 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 126 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 126 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 125.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 125.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 125.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 125.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 125.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 125.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 125.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 125.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 125.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 125.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 125.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 125.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 125.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 125.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 125.616 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 125.426 13.39 126.574 ;
      VIA 12.576 126.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 126.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 126.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 126.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 126.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 126.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 126.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 126.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 126.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 126.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 126.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 126.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 126.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 126.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 126.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 126 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 126 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 126 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 126 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 126 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 125.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 125.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 125.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 125.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 125.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 125.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 125.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 125.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 125.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 125.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 125.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 125.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 125.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 125.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 125.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 126 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 116.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 116.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 116.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 116.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 116.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 116.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 116.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 116.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 116.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 116.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 116.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 116.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 116.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 116.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 116.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 115.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 115.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 115.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 115.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 115.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 115.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 115.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 115.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 115.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 115.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 115.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 115.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 115.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 115.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 115.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 115.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 115.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 115.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 115.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 115.536 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 115.346 13.39 116.494 ;
      VIA 12.576 116.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 116.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 116.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 116.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 116.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 116.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 116.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 116.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 116.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 116.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 116.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 116.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 116.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 116.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 116.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 115.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 115.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 115.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 115.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 115.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 115.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 115.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 115.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 115.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 115.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 115.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 115.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 115.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 115.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 115.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 115.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 115.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 115.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 115.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 115.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 115.92 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 106.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 106.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 106.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 106.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 106.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 106.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 106.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 106.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 106.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 106.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 105.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 105.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 105.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 105.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 105.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 105.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 105.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 105.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 105.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 105.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 105.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 105.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 105.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 105.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 105.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 105.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 105.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 105.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 105.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 105.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 105.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 105.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 105.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 105.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 105.456 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 105.266 13.39 106.414 ;
      VIA 12.576 106.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 106.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 106.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 106.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 106.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 106.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 106.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 106.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 106.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 106.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 105.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 105.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 105.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 105.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 105.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 105.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 105.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 105.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 105.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 105.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 105.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 105.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 105.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 105.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 105.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 105.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 105.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 105.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 105.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 105.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 105.84 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 96.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 96.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 96.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 96.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 96.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 96.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 96.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 96.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 96.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 96.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 95.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 95.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 95.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 95.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 95.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 95.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 95.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 95.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 95.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 95.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 95.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 95.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 95.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 95.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 95.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 95.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 95.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 95.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 95.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 95.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 95.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 95.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 95.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 95.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 95.376 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 95.186 13.39 96.334 ;
      VIA 12.576 96.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 96.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 96.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 96.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 96.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 96.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 96.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 96.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 96.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 96.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 95.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 95.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 95.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 95.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 95.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 95.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 95.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 95.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 95.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 95.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 95.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 95.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 95.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 95.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 95.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 95.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 95.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 95.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 95.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 95.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 95.76 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 86.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 86.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 86.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 86.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 86.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 85.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 85.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 85.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 85.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 85.296 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 85.106 13.39 86.254 ;
      VIA 12.576 86.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 86.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 86.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 86.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 86.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 85.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 85.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 85.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 85.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 85.68 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 75.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 75.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 75.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 75.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 75.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 75.216 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 75.026 13.39 76.174 ;
      VIA 12.576 75.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 75.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 75.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 75.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 75.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 75.6 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 65.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 65.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 65.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 65.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 65.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 65.136 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 64.946 13.39 66.094 ;
      VIA 12.576 65.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 65.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 65.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 65.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 65.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 65.52 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 55.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 55.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 55.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 55.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 55.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 55.056 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 54.866 13.39 56.014 ;
      VIA 12.576 55.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 55.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 55.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 55.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 55.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 55.44 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 45.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 45.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 45.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 45.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 45.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 45.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 45.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 45.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 45.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 45.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 44.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 44.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 44.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 44.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 44.976 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 44.786 13.39 45.934 ;
      VIA 12.576 45.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 45.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 45.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 45.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 45.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 45.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 45.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 45.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 45.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 44.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 44.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 44.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 44.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 44.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 45.36 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 35.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 35.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 35.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 35.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 35.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 35.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 35.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 35.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 35.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 35.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 34.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 34.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 34.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 34.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 34.896 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 34.706 13.39 35.854 ;
      VIA 12.576 35.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 35.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 35.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 35.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 35.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 35.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 35.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 35.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 35.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 34.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 34.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 34.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 34.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 34.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 35.28 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 25.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 25.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 25.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 25.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 25.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 25.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 25.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 25.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 25.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 25.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 25.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 25.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 25.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 25.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 25.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 25.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 25.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 25.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 25.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 25.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 25.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 25.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 25.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 25.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 25.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 24.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 24.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 24.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 24.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 24.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 24.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 24.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 24.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 24.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 24.816 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 24.626 13.39 25.774 ;
      VIA 12.576 25.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 25.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 25.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 25.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 25.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 25.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 25.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 25.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 25.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 25.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 25.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 25.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 25.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 25.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 25.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 25.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 25.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 25.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 25.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 25.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 24.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 24.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 24.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 24.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 24.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 24.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 24.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 24.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 24.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 24.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 25.2 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 12.856 15.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 15.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 15.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 15.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 15.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 15.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 15.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 15.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 15.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 15.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 15.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 15.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 15.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 15.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 15.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 15.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 15.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 15.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 15.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 15.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 14.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 14.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 14.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 14.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 14.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 14.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 14.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 14.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 14.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 14.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.856 14.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.728 14.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.6 14.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.472 14.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 12.344 14.736 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  11.25 14.546 13.39 15.694 ;
      VIA 12.576 15.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 15.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 15.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 15.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 15.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 15.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 15.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 15.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 15.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 15.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 15.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 15.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 15.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 15.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 15.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 15.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 15.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 15.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 15.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 15.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 14.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 14.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 14.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 14.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 14.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 14.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 14.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 14.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 14.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 14.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.576 14.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.448 14.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 14.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.192 14.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.064 14.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 12.32 15.12 via1_2_4480_1800_1_4_1240_1240 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  997.66 9.506 1002.14 262.654 ;
        RECT  14.18 342.146 16.42 595.294 ;
        RECT  997.66 342.146 1002.14 595.294 ;
        RECT  14.18 9.506 16.42 262.654 ;
        RECT  971.04 9.506 975.52 605.374 ;
        RECT  926.24 9.506 930.72 605.374 ;
        RECT  881.44 9.506 885.92 605.374 ;
        RECT  836.64 9.506 841.12 605.374 ;
        RECT  791.84 9.506 796.32 605.374 ;
        RECT  747.04 9.506 751.52 605.374 ;
        RECT  702.24 9.506 706.72 605.374 ;
        RECT  657.44 9.506 661.92 605.374 ;
        RECT  612.64 9.506 617.12 605.374 ;
        RECT  567.84 9.506 572.32 605.374 ;
        RECT  523.04 9.506 527.52 605.374 ;
        RECT  478.24 9.506 482.72 605.374 ;
        RECT  433.44 9.506 437.92 605.374 ;
        RECT  388.64 9.506 393.12 605.374 ;
        RECT  343.84 9.506 348.32 605.374 ;
        RECT  299.04 9.506 303.52 605.374 ;
        RECT  254.24 9.506 258.72 605.374 ;
        RECT  209.44 9.506 213.92 605.374 ;
        RECT  164.64 9.506 169.12 605.374 ;
        RECT  119.84 9.506 124.32 605.374 ;
        RECT  75.04 9.506 79.52 605.374 ;
        RECT  30.24 9.506 34.72 605.374 ;
      LAYER Metal1 ;
        RECT  985.04 584.19 1009.68 585.09 ;
        RECT  985.04 574.11 1009.68 575.01 ;
        RECT  985.04 564.03 1009.68 564.93 ;
        RECT  985.04 553.95 1009.68 554.85 ;
        RECT  985.04 543.87 1009.68 544.77 ;
        RECT  985.04 533.79 1009.68 534.69 ;
        RECT  985.04 523.71 1009.68 524.61 ;
        RECT  985.04 513.63 1009.68 514.53 ;
        RECT  985.04 503.55 1009.68 504.45 ;
        RECT  985.04 493.47 1009.68 494.37 ;
        RECT  985.04 483.39 1009.68 484.29 ;
        RECT  985.04 473.31 1009.68 474.21 ;
        RECT  985.04 463.23 1009.68 464.13 ;
        RECT  985.04 453.15 1009.68 454.05 ;
        RECT  985.04 443.07 1009.68 443.97 ;
        RECT  985.04 432.99 1009.68 433.89 ;
        RECT  985.04 422.91 1009.68 423.81 ;
        RECT  985.04 412.83 1009.68 413.73 ;
        RECT  985.04 402.75 1009.68 403.65 ;
        RECT  985.04 392.67 1009.68 393.57 ;
        RECT  985.04 382.59 1009.68 383.49 ;
        RECT  985.04 372.51 1009.68 373.41 ;
        RECT  985.04 362.43 1009.68 363.33 ;
        RECT  985.04 352.35 1009.68 353.25 ;
        RECT  985.04 251.55 1009.68 252.45 ;
        RECT  985.04 241.47 1009.68 242.37 ;
        RECT  985.04 231.39 1009.68 232.29 ;
        RECT  985.04 221.31 1009.68 222.21 ;
        RECT  985.04 211.23 1009.68 212.13 ;
        RECT  985.04 201.15 1009.68 202.05 ;
        RECT  985.04 191.07 1009.68 191.97 ;
        RECT  985.04 180.99 1009.68 181.89 ;
        RECT  985.04 170.91 1009.68 171.81 ;
        RECT  985.04 160.83 1009.68 161.73 ;
        RECT  985.04 150.75 1009.68 151.65 ;
        RECT  985.04 140.67 1009.68 141.57 ;
        RECT  985.04 130.59 1009.68 131.49 ;
        RECT  985.04 120.51 1009.68 121.41 ;
        RECT  985.04 110.43 1009.68 111.33 ;
        RECT  985.04 100.35 1009.68 101.25 ;
        RECT  985.04 90.27 1009.68 91.17 ;
        RECT  985.04 80.19 1009.68 81.09 ;
        RECT  985.04 70.11 1009.68 71.01 ;
        RECT  985.04 60.03 1009.68 60.93 ;
        RECT  985.04 49.95 1009.68 50.85 ;
        RECT  985.04 39.87 1009.68 40.77 ;
        RECT  985.04 29.79 1009.68 30.69 ;
        RECT  985.04 19.71 1009.68 20.61 ;
        RECT  454.16 584.19 548.8 585.09 ;
        RECT  454.16 574.11 548.8 575.01 ;
        RECT  454.16 564.03 548.8 564.93 ;
        RECT  454.16 553.95 548.8 554.85 ;
        RECT  454.16 543.87 548.8 544.77 ;
        RECT  454.16 533.79 548.8 534.69 ;
        RECT  454.16 523.71 548.8 524.61 ;
        RECT  454.16 513.63 548.8 514.53 ;
        RECT  454.16 503.55 548.8 504.45 ;
        RECT  454.16 493.47 548.8 494.37 ;
        RECT  454.16 483.39 548.8 484.29 ;
        RECT  454.16 473.31 548.8 474.21 ;
        RECT  454.16 463.23 548.8 464.13 ;
        RECT  454.16 453.15 548.8 454.05 ;
        RECT  454.16 443.07 548.8 443.97 ;
        RECT  454.16 432.99 548.8 433.89 ;
        RECT  454.16 422.91 548.8 423.81 ;
        RECT  454.16 412.83 548.8 413.73 ;
        RECT  454.16 402.75 548.8 403.65 ;
        RECT  454.16 392.67 548.8 393.57 ;
        RECT  454.16 382.59 548.8 383.49 ;
        RECT  454.16 372.51 548.8 373.41 ;
        RECT  454.16 362.43 548.8 363.33 ;
        RECT  454.16 352.35 548.8 353.25 ;
        RECT  454.16 251.55 548.8 252.45 ;
        RECT  454.16 241.47 548.8 242.37 ;
        RECT  454.16 231.39 548.8 232.29 ;
        RECT  454.16 221.31 548.8 222.21 ;
        RECT  454.16 211.23 548.8 212.13 ;
        RECT  454.16 201.15 548.8 202.05 ;
        RECT  454.16 191.07 548.8 191.97 ;
        RECT  454.16 180.99 548.8 181.89 ;
        RECT  454.16 170.91 548.8 171.81 ;
        RECT  454.16 160.83 548.8 161.73 ;
        RECT  454.16 150.75 548.8 151.65 ;
        RECT  454.16 140.67 548.8 141.57 ;
        RECT  454.16 130.59 548.8 131.49 ;
        RECT  454.16 120.51 548.8 121.41 ;
        RECT  454.16 110.43 548.8 111.33 ;
        RECT  454.16 100.35 548.8 101.25 ;
        RECT  454.16 90.27 548.8 91.17 ;
        RECT  454.16 80.19 548.8 81.09 ;
        RECT  454.16 70.11 548.8 71.01 ;
        RECT  454.16 60.03 548.8 60.93 ;
        RECT  454.16 49.95 548.8 50.85 ;
        RECT  454.16 39.87 548.8 40.77 ;
        RECT  454.16 29.79 548.8 30.69 ;
        RECT  454.16 19.71 548.8 20.61 ;
        RECT  10.08 604.35 1009.68 605.25 ;
        RECT  10.08 594.27 1009.68 595.17 ;
        RECT  10.08 584.19 17.92 585.09 ;
        RECT  10.08 574.11 17.92 575.01 ;
        RECT  10.08 564.03 17.92 564.93 ;
        RECT  10.08 553.95 17.92 554.85 ;
        RECT  10.08 543.87 17.92 544.77 ;
        RECT  10.08 533.79 17.92 534.69 ;
        RECT  10.08 523.71 17.92 524.61 ;
        RECT  10.08 513.63 17.92 514.53 ;
        RECT  10.08 503.55 17.92 504.45 ;
        RECT  10.08 493.47 17.92 494.37 ;
        RECT  10.08 483.39 17.92 484.29 ;
        RECT  10.08 473.31 17.92 474.21 ;
        RECT  10.08 463.23 17.92 464.13 ;
        RECT  10.08 453.15 17.92 454.05 ;
        RECT  10.08 443.07 17.92 443.97 ;
        RECT  10.08 432.99 17.92 433.89 ;
        RECT  10.08 422.91 17.92 423.81 ;
        RECT  10.08 412.83 17.92 413.73 ;
        RECT  10.08 402.75 17.92 403.65 ;
        RECT  10.08 392.67 17.92 393.57 ;
        RECT  10.08 382.59 17.92 383.49 ;
        RECT  10.08 372.51 17.92 373.41 ;
        RECT  10.08 362.43 17.92 363.33 ;
        RECT  10.08 352.35 17.92 353.25 ;
        RECT  10.08 342.27 1009.68 343.17 ;
        RECT  10.08 332.19 1009.68 333.09 ;
        RECT  10.08 322.11 1009.68 323.01 ;
        RECT  10.08 312.03 1009.68 312.93 ;
        RECT  10.08 301.95 1009.68 302.85 ;
        RECT  10.08 291.87 1009.68 292.77 ;
        RECT  10.08 281.79 1009.68 282.69 ;
        RECT  10.08 271.71 1009.68 272.61 ;
        RECT  10.08 261.63 1009.68 262.53 ;
        RECT  10.08 251.55 17.92 252.45 ;
        RECT  10.08 241.47 17.92 242.37 ;
        RECT  10.08 231.39 17.92 232.29 ;
        RECT  10.08 221.31 17.92 222.21 ;
        RECT  10.08 211.23 17.92 212.13 ;
        RECT  10.08 201.15 17.92 202.05 ;
        RECT  10.08 191.07 17.92 191.97 ;
        RECT  10.08 180.99 17.92 181.89 ;
        RECT  10.08 170.91 17.92 171.81 ;
        RECT  10.08 160.83 17.92 161.73 ;
        RECT  10.08 150.75 17.92 151.65 ;
        RECT  10.08 140.67 17.92 141.57 ;
        RECT  10.08 130.59 17.92 131.49 ;
        RECT  10.08 120.51 17.92 121.41 ;
        RECT  10.08 110.43 17.92 111.33 ;
        RECT  10.08 100.35 17.92 101.25 ;
        RECT  10.08 90.27 17.92 91.17 ;
        RECT  10.08 80.19 17.92 81.09 ;
        RECT  10.08 70.11 17.92 71.01 ;
        RECT  10.08 60.03 17.92 60.93 ;
        RECT  10.08 49.95 17.92 50.85 ;
        RECT  10.08 39.87 17.92 40.77 ;
        RECT  10.08 29.79 17.92 30.69 ;
        RECT  10.08 19.71 17.92 20.61 ;
        RECT  10.08 9.63 1009.68 10.53 ;
      VIA 1000.156 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 594.146 1001.23 595.294 ;
      VIA 1000.416 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 584.066 1001.23 585.214 ;
      VIA 1000.416 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 573.986 1001.23 575.134 ;
      VIA 1000.416 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 563.906 1001.23 565.054 ;
      VIA 1000.416 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 553.826 1001.23 554.974 ;
      VIA 1000.416 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 543.746 1001.23 544.894 ;
      VIA 1000.416 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 533.666 1001.23 534.814 ;
      VIA 1000.416 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 523.586 1001.23 524.734 ;
      VIA 1000.416 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 513.506 1001.23 514.654 ;
      VIA 1000.416 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 503.426 1001.23 504.574 ;
      VIA 1000.416 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 493.346 1001.23 494.494 ;
      VIA 1000.416 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 483.266 1001.23 484.414 ;
      VIA 1000.416 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 473.186 1001.23 474.334 ;
      VIA 1000.416 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 463.106 1001.23 464.254 ;
      VIA 1000.416 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 453.026 1001.23 454.174 ;
      VIA 1000.416 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 442.946 1001.23 444.094 ;
      VIA 1000.416 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 432.866 1001.23 434.014 ;
      VIA 1000.416 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 422.786 1001.23 423.934 ;
      VIA 1000.416 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 412.706 1001.23 413.854 ;
      VIA 1000.416 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 402.626 1001.23 403.774 ;
      VIA 1000.416 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 392.546 1001.23 393.694 ;
      VIA 1000.416 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 382.466 1001.23 383.614 ;
      VIA 1000.416 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 372.386 1001.23 373.534 ;
      VIA 1000.416 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 362.306 1001.23 363.454 ;
      VIA 1000.416 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 352.226 1001.23 353.374 ;
      VIA 1000.416 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 342.146 1001.23 343.294 ;
      VIA 1000.416 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 261.506 1001.23 262.654 ;
      VIA 1000.416 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 251.426 1001.23 252.574 ;
      VIA 1000.416 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 241.346 1001.23 242.494 ;
      VIA 1000.416 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 231.266 1001.23 232.414 ;
      VIA 1000.416 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 221.186 1001.23 222.334 ;
      VIA 1000.416 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 211.106 1001.23 212.254 ;
      VIA 1000.416 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 201.026 1001.23 202.174 ;
      VIA 1000.416 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 190.946 1001.23 192.094 ;
      VIA 1000.416 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 180.866 1001.23 182.014 ;
      VIA 1000.416 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 170.786 1001.23 171.934 ;
      VIA 1000.416 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 160.706 1001.23 161.854 ;
      VIA 1000.416 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 150.626 1001.23 151.774 ;
      VIA 1000.416 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 140.546 1001.23 141.694 ;
      VIA 1000.416 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 130.466 1001.23 131.614 ;
      VIA 1000.416 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 120.386 1001.23 121.534 ;
      VIA 1000.416 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 110.306 1001.23 111.454 ;
      VIA 1000.416 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 100.226 1001.23 101.374 ;
      VIA 1000.416 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 90.146 1001.23 91.294 ;
      VIA 1000.416 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 80.066 1001.23 81.214 ;
      VIA 1000.416 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 69.986 1001.23 71.134 ;
      VIA 1000.416 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 59.906 1001.23 61.054 ;
      VIA 1000.416 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 49.826 1001.23 50.974 ;
      VIA 1000.416 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 39.746 1001.23 40.894 ;
      VIA 1000.416 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 29.666 1001.23 30.814 ;
      VIA 1000.416 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 19.586 1001.23 20.734 ;
      VIA 1000.416 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 1000.156 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.156 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 1000.028 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.9 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.772 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 999.644 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  999.09 9.506 1001.23 10.654 ;
      VIA 1000.416 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.416 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.288 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.032 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 999.904 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 1000.16 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 604.226 974.35 605.374 ;
      VIA 973.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 594.146 974.35 595.294 ;
      VIA 973.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 342.146 974.35 343.294 ;
      VIA 973.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 332.066 974.35 333.214 ;
      VIA 973.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 321.986 974.35 323.134 ;
      VIA 973.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 311.906 974.35 313.054 ;
      VIA 973.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 301.826 974.35 302.974 ;
      VIA 973.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 291.746 974.35 292.894 ;
      VIA 973.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 281.666 974.35 282.814 ;
      VIA 973.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 271.586 974.35 272.734 ;
      VIA 973.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 261.506 974.35 262.654 ;
      VIA 973.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 973.156 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.156 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 973.028 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.9 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.772 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 972.644 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  972.21 9.506 974.35 10.654 ;
      VIA 973.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 973.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 604.226 929.55 605.374 ;
      VIA 928.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 594.146 929.55 595.294 ;
      VIA 928.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 342.146 929.55 343.294 ;
      VIA 928.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 332.066 929.55 333.214 ;
      VIA 928.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 321.986 929.55 323.134 ;
      VIA 928.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 311.906 929.55 313.054 ;
      VIA 928.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 301.826 929.55 302.974 ;
      VIA 928.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 291.746 929.55 292.894 ;
      VIA 928.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 281.666 929.55 282.814 ;
      VIA 928.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 271.586 929.55 272.734 ;
      VIA 928.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 261.506 929.55 262.654 ;
      VIA 928.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 929.056 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 929.056 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.928 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.8 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.672 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 928.544 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  927.41 9.506 929.55 10.654 ;
      VIA 928.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 928.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 604.226 884.75 605.374 ;
      VIA 883.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 594.146 884.75 595.294 ;
      VIA 883.936 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 342.146 884.75 343.294 ;
      VIA 883.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 332.066 884.75 333.214 ;
      VIA 883.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 321.986 884.75 323.134 ;
      VIA 883.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 311.906 884.75 313.054 ;
      VIA 883.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 301.826 884.75 302.974 ;
      VIA 883.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 291.746 884.75 292.894 ;
      VIA 883.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 281.666 884.75 282.814 ;
      VIA 883.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 271.586 884.75 272.734 ;
      VIA 883.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 261.506 884.75 262.654 ;
      VIA 883.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 884.056 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 884.056 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.928 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.8 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.672 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 883.544 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  882.61 9.506 884.75 10.654 ;
      VIA 883.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 883.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 604.226 839.95 605.374 ;
      VIA 839.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 594.146 839.95 595.294 ;
      VIA 839.136 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 342.146 839.95 343.294 ;
      VIA 839.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 332.066 839.95 333.214 ;
      VIA 839.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 321.986 839.95 323.134 ;
      VIA 839.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 311.906 839.95 313.054 ;
      VIA 839.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 301.826 839.95 302.974 ;
      VIA 839.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 291.746 839.95 292.894 ;
      VIA 839.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 281.666 839.95 282.814 ;
      VIA 839.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 271.586 839.95 272.734 ;
      VIA 839.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 261.506 839.95 262.654 ;
      VIA 839.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 839.056 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 839.056 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.928 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.8 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.672 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 838.544 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  837.81 9.506 839.95 10.654 ;
      VIA 839.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 839.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 838.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 604.226 795.15 605.374 ;
      VIA 794.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 594.146 795.15 595.294 ;
      VIA 794.336 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 342.146 795.15 343.294 ;
      VIA 794.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 332.066 795.15 333.214 ;
      VIA 794.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 321.986 795.15 323.134 ;
      VIA 794.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 311.906 795.15 313.054 ;
      VIA 794.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 301.826 795.15 302.974 ;
      VIA 794.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 291.746 795.15 292.894 ;
      VIA 794.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 281.666 795.15 282.814 ;
      VIA 794.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 271.586 795.15 272.734 ;
      VIA 794.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 261.506 795.15 262.654 ;
      VIA 794.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 794.056 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 794.056 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.928 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.8 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.672 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 793.544 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  793.01 9.506 795.15 10.654 ;
      VIA 794.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 793.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 794.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 604.226 750.35 605.374 ;
      VIA 749.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 594.146 750.35 595.294 ;
      VIA 749.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 342.146 750.35 343.294 ;
      VIA 749.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 332.066 750.35 333.214 ;
      VIA 749.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 321.986 750.35 323.134 ;
      VIA 749.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 311.906 750.35 313.054 ;
      VIA 749.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 301.826 750.35 302.974 ;
      VIA 749.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 291.746 750.35 292.894 ;
      VIA 749.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 281.666 750.35 282.814 ;
      VIA 749.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 271.586 750.35 272.734 ;
      VIA 749.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 261.506 750.35 262.654 ;
      VIA 749.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 749.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 749.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  748.21 9.506 750.35 10.654 ;
      VIA 749.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 749.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 604.226 705.55 605.374 ;
      VIA 704.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 594.146 705.55 595.294 ;
      VIA 704.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 342.146 705.55 343.294 ;
      VIA 704.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 332.066 705.55 333.214 ;
      VIA 704.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 321.986 705.55 323.134 ;
      VIA 704.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 311.906 705.55 313.054 ;
      VIA 704.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 301.826 705.55 302.974 ;
      VIA 704.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 291.746 705.55 292.894 ;
      VIA 704.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 281.666 705.55 282.814 ;
      VIA 704.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 271.586 705.55 272.734 ;
      VIA 704.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 261.506 705.55 262.654 ;
      VIA 704.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 704.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 704.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  703.41 9.506 705.55 10.654 ;
      VIA 704.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 704.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 604.226 660.75 605.374 ;
      VIA 659.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 594.146 660.75 595.294 ;
      VIA 659.936 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 342.146 660.75 343.294 ;
      VIA 659.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 332.066 660.75 333.214 ;
      VIA 659.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 321.986 660.75 323.134 ;
      VIA 659.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 311.906 660.75 313.054 ;
      VIA 659.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 301.826 660.75 302.974 ;
      VIA 659.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 291.746 660.75 292.894 ;
      VIA 659.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 281.666 660.75 282.814 ;
      VIA 659.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 271.586 660.75 272.734 ;
      VIA 659.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 261.506 660.75 262.654 ;
      VIA 659.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 659.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 659.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  658.61 9.506 660.75 10.654 ;
      VIA 659.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 659.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 604.226 615.95 605.374 ;
      VIA 615.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 594.146 615.95 595.294 ;
      VIA 615.136 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 342.146 615.95 343.294 ;
      VIA 615.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 332.066 615.95 333.214 ;
      VIA 615.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 321.986 615.95 323.134 ;
      VIA 615.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 311.906 615.95 313.054 ;
      VIA 615.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 301.826 615.95 302.974 ;
      VIA 615.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 291.746 615.95 292.894 ;
      VIA 615.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 281.666 615.95 282.814 ;
      VIA 615.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 271.586 615.95 272.734 ;
      VIA 615.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 261.506 615.95 262.654 ;
      VIA 615.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 614.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 614.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  613.81 9.506 615.95 10.654 ;
      VIA 615.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 615.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 614.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 604.226 571.15 605.374 ;
      VIA 570.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 594.146 571.15 595.294 ;
      VIA 570.336 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 342.146 571.15 343.294 ;
      VIA 570.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 332.066 571.15 333.214 ;
      VIA 570.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 321.986 571.15 323.134 ;
      VIA 570.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 311.906 571.15 313.054 ;
      VIA 570.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 301.826 571.15 302.974 ;
      VIA 570.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 291.746 571.15 292.894 ;
      VIA 570.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 281.666 571.15 282.814 ;
      VIA 570.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 271.586 571.15 272.734 ;
      VIA 570.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 261.506 571.15 262.654 ;
      VIA 570.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 9.506 571.15 10.654 ;
      VIA 570.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 604.226 526.35 605.374 ;
      VIA 525.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 594.146 526.35 595.294 ;
      VIA 525.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 584.066 526.35 585.214 ;
      VIA 525.536 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 573.986 526.35 575.134 ;
      VIA 525.536 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 563.906 526.35 565.054 ;
      VIA 525.536 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 553.826 526.35 554.974 ;
      VIA 525.536 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 543.746 526.35 544.894 ;
      VIA 525.536 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 533.666 526.35 534.814 ;
      VIA 525.536 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 523.586 526.35 524.734 ;
      VIA 525.536 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 513.506 526.35 514.654 ;
      VIA 525.536 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 503.426 526.35 504.574 ;
      VIA 525.536 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 493.346 526.35 494.494 ;
      VIA 525.536 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 483.266 526.35 484.414 ;
      VIA 525.536 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 473.186 526.35 474.334 ;
      VIA 525.536 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 463.106 526.35 464.254 ;
      VIA 525.536 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 453.026 526.35 454.174 ;
      VIA 525.536 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 442.946 526.35 444.094 ;
      VIA 525.536 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 432.866 526.35 434.014 ;
      VIA 525.536 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 422.786 526.35 423.934 ;
      VIA 525.536 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 412.706 526.35 413.854 ;
      VIA 525.536 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 402.626 526.35 403.774 ;
      VIA 525.536 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 392.546 526.35 393.694 ;
      VIA 525.536 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 382.466 526.35 383.614 ;
      VIA 525.536 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 372.386 526.35 373.534 ;
      VIA 525.536 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 362.306 526.35 363.454 ;
      VIA 525.536 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 352.226 526.35 353.374 ;
      VIA 525.536 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 342.146 526.35 343.294 ;
      VIA 525.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 332.066 526.35 333.214 ;
      VIA 525.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 321.986 526.35 323.134 ;
      VIA 525.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 311.906 526.35 313.054 ;
      VIA 525.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 301.826 526.35 302.974 ;
      VIA 525.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 291.746 526.35 292.894 ;
      VIA 525.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 281.666 526.35 282.814 ;
      VIA 525.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 271.586 526.35 272.734 ;
      VIA 525.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 261.506 526.35 262.654 ;
      VIA 525.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 251.426 526.35 252.574 ;
      VIA 525.536 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 241.346 526.35 242.494 ;
      VIA 525.536 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 231.266 526.35 232.414 ;
      VIA 525.536 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 221.186 526.35 222.334 ;
      VIA 525.536 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 211.106 526.35 212.254 ;
      VIA 525.536 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 201.026 526.35 202.174 ;
      VIA 525.536 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 190.946 526.35 192.094 ;
      VIA 525.536 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 180.866 526.35 182.014 ;
      VIA 525.536 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 170.786 526.35 171.934 ;
      VIA 525.536 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 160.706 526.35 161.854 ;
      VIA 525.536 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 150.626 526.35 151.774 ;
      VIA 525.536 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 140.546 526.35 141.694 ;
      VIA 525.536 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 130.466 526.35 131.614 ;
      VIA 525.536 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 120.386 526.35 121.534 ;
      VIA 525.536 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 110.306 526.35 111.454 ;
      VIA 525.536 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 100.226 526.35 101.374 ;
      VIA 525.536 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 90.146 526.35 91.294 ;
      VIA 525.536 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 80.066 526.35 81.214 ;
      VIA 525.536 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 69.986 526.35 71.134 ;
      VIA 525.536 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 59.906 526.35 61.054 ;
      VIA 525.536 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 49.826 526.35 50.974 ;
      VIA 525.536 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 39.746 526.35 40.894 ;
      VIA 525.536 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 29.666 526.35 30.814 ;
      VIA 525.536 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 19.586 526.35 20.734 ;
      VIA 525.536 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 9.506 526.35 10.654 ;
      VIA 525.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 604.226 481.55 605.374 ;
      VIA 480.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 594.146 481.55 595.294 ;
      VIA 480.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 584.066 481.55 585.214 ;
      VIA 480.736 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 573.986 481.55 575.134 ;
      VIA 480.736 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 563.906 481.55 565.054 ;
      VIA 480.736 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 553.826 481.55 554.974 ;
      VIA 480.736 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 543.746 481.55 544.894 ;
      VIA 480.736 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 533.666 481.55 534.814 ;
      VIA 480.736 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 523.586 481.55 524.734 ;
      VIA 480.736 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 513.506 481.55 514.654 ;
      VIA 480.736 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 503.426 481.55 504.574 ;
      VIA 480.736 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 493.346 481.55 494.494 ;
      VIA 480.736 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 483.266 481.55 484.414 ;
      VIA 480.736 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 473.186 481.55 474.334 ;
      VIA 480.736 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 463.106 481.55 464.254 ;
      VIA 480.736 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 453.026 481.55 454.174 ;
      VIA 480.736 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 442.946 481.55 444.094 ;
      VIA 480.736 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 432.866 481.55 434.014 ;
      VIA 480.736 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 422.786 481.55 423.934 ;
      VIA 480.736 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 412.706 481.55 413.854 ;
      VIA 480.736 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 402.626 481.55 403.774 ;
      VIA 480.736 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 392.546 481.55 393.694 ;
      VIA 480.736 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 382.466 481.55 383.614 ;
      VIA 480.736 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 372.386 481.55 373.534 ;
      VIA 480.736 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 362.306 481.55 363.454 ;
      VIA 480.736 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 352.226 481.55 353.374 ;
      VIA 480.736 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 342.146 481.55 343.294 ;
      VIA 480.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 332.066 481.55 333.214 ;
      VIA 480.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 321.986 481.55 323.134 ;
      VIA 480.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 311.906 481.55 313.054 ;
      VIA 480.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 301.826 481.55 302.974 ;
      VIA 480.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 291.746 481.55 292.894 ;
      VIA 480.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 281.666 481.55 282.814 ;
      VIA 480.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 271.586 481.55 272.734 ;
      VIA 480.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 261.506 481.55 262.654 ;
      VIA 480.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 251.426 481.55 252.574 ;
      VIA 480.736 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 241.346 481.55 242.494 ;
      VIA 480.736 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 231.266 481.55 232.414 ;
      VIA 480.736 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 221.186 481.55 222.334 ;
      VIA 480.736 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 211.106 481.55 212.254 ;
      VIA 480.736 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 201.026 481.55 202.174 ;
      VIA 480.736 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 190.946 481.55 192.094 ;
      VIA 480.736 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 180.866 481.55 182.014 ;
      VIA 480.736 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 170.786 481.55 171.934 ;
      VIA 480.736 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 160.706 481.55 161.854 ;
      VIA 480.736 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 150.626 481.55 151.774 ;
      VIA 480.736 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 140.546 481.55 141.694 ;
      VIA 480.736 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 130.466 481.55 131.614 ;
      VIA 480.736 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 120.386 481.55 121.534 ;
      VIA 480.736 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 110.306 481.55 111.454 ;
      VIA 480.736 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 100.226 481.55 101.374 ;
      VIA 480.736 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 90.146 481.55 91.294 ;
      VIA 480.736 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 80.066 481.55 81.214 ;
      VIA 480.736 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 69.986 481.55 71.134 ;
      VIA 480.736 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 59.906 481.55 61.054 ;
      VIA 480.736 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 49.826 481.55 50.974 ;
      VIA 480.736 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 39.746 481.55 40.894 ;
      VIA 480.736 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 29.666 481.55 30.814 ;
      VIA 480.736 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 19.586 481.55 20.734 ;
      VIA 480.736 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 9.506 481.55 10.654 ;
      VIA 480.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 604.226 436.75 605.374 ;
      VIA 435.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 594.146 436.75 595.294 ;
      VIA 435.936 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 342.146 436.75 343.294 ;
      VIA 435.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 332.066 436.75 333.214 ;
      VIA 435.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 321.986 436.75 323.134 ;
      VIA 435.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 311.906 436.75 313.054 ;
      VIA 435.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 301.826 436.75 302.974 ;
      VIA 435.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 291.746 436.75 292.894 ;
      VIA 435.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 281.666 436.75 282.814 ;
      VIA 435.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 271.586 436.75 272.734 ;
      VIA 435.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 261.506 436.75 262.654 ;
      VIA 435.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 9.506 436.75 10.654 ;
      VIA 435.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 604.226 391.95 605.374 ;
      VIA 391.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 594.146 391.95 595.294 ;
      VIA 391.136 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 342.146 391.95 343.294 ;
      VIA 391.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 332.066 391.95 333.214 ;
      VIA 391.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 321.986 391.95 323.134 ;
      VIA 391.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 311.906 391.95 313.054 ;
      VIA 391.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 301.826 391.95 302.974 ;
      VIA 391.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 291.746 391.95 292.894 ;
      VIA 391.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 281.666 391.95 282.814 ;
      VIA 391.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 271.586 391.95 272.734 ;
      VIA 391.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 261.506 391.95 262.654 ;
      VIA 391.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 9.506 391.95 10.654 ;
      VIA 391.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 604.226 347.15 605.374 ;
      VIA 346.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 594.146 347.15 595.294 ;
      VIA 346.336 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 342.146 347.15 343.294 ;
      VIA 346.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 332.066 347.15 333.214 ;
      VIA 346.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 321.986 347.15 323.134 ;
      VIA 346.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 311.906 347.15 313.054 ;
      VIA 346.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 301.826 347.15 302.974 ;
      VIA 346.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 291.746 347.15 292.894 ;
      VIA 346.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 281.666 347.15 282.814 ;
      VIA 346.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 271.586 347.15 272.734 ;
      VIA 346.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 261.506 347.15 262.654 ;
      VIA 346.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 9.506 347.15 10.654 ;
      VIA 346.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 604.226 302.35 605.374 ;
      VIA 301.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 594.146 302.35 595.294 ;
      VIA 301.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 342.146 302.35 343.294 ;
      VIA 301.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 332.066 302.35 333.214 ;
      VIA 301.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 321.986 302.35 323.134 ;
      VIA 301.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 311.906 302.35 313.054 ;
      VIA 301.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 301.826 302.35 302.974 ;
      VIA 301.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 291.746 302.35 292.894 ;
      VIA 301.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 281.666 302.35 282.814 ;
      VIA 301.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 271.586 302.35 272.734 ;
      VIA 301.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 261.506 302.35 262.654 ;
      VIA 301.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 9.506 302.35 10.654 ;
      VIA 301.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 604.226 257.55 605.374 ;
      VIA 256.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 594.146 257.55 595.294 ;
      VIA 256.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 342.146 257.55 343.294 ;
      VIA 256.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 332.066 257.55 333.214 ;
      VIA 256.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 321.986 257.55 323.134 ;
      VIA 256.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 311.906 257.55 313.054 ;
      VIA 256.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 301.826 257.55 302.974 ;
      VIA 256.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 291.746 257.55 292.894 ;
      VIA 256.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 281.666 257.55 282.814 ;
      VIA 256.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 271.586 257.55 272.734 ;
      VIA 256.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 261.506 257.55 262.654 ;
      VIA 256.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 9.506 257.55 10.654 ;
      VIA 256.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 604.226 212.75 605.374 ;
      VIA 211.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 594.146 212.75 595.294 ;
      VIA 211.936 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 342.146 212.75 343.294 ;
      VIA 211.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 332.066 212.75 333.214 ;
      VIA 211.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 321.986 212.75 323.134 ;
      VIA 211.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 311.906 212.75 313.054 ;
      VIA 211.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 301.826 212.75 302.974 ;
      VIA 211.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 291.746 212.75 292.894 ;
      VIA 211.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 281.666 212.75 282.814 ;
      VIA 211.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 271.586 212.75 272.734 ;
      VIA 211.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 261.506 212.75 262.654 ;
      VIA 211.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 9.506 212.75 10.654 ;
      VIA 211.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 604.226 167.95 605.374 ;
      VIA 167.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 594.146 167.95 595.294 ;
      VIA 167.136 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 342.146 167.95 343.294 ;
      VIA 167.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 332.066 167.95 333.214 ;
      VIA 167.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 321.986 167.95 323.134 ;
      VIA 167.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 311.906 167.95 313.054 ;
      VIA 167.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 301.826 167.95 302.974 ;
      VIA 167.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 291.746 167.95 292.894 ;
      VIA 167.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 281.666 167.95 282.814 ;
      VIA 167.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 271.586 167.95 272.734 ;
      VIA 167.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 261.506 167.95 262.654 ;
      VIA 167.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 9.506 167.95 10.654 ;
      VIA 167.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 604.226 123.15 605.374 ;
      VIA 122.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 594.146 123.15 595.294 ;
      VIA 122.336 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 342.146 123.15 343.294 ;
      VIA 122.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 332.066 123.15 333.214 ;
      VIA 122.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 321.986 123.15 323.134 ;
      VIA 122.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 311.906 123.15 313.054 ;
      VIA 122.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 301.826 123.15 302.974 ;
      VIA 122.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 291.746 123.15 292.894 ;
      VIA 122.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 281.666 123.15 282.814 ;
      VIA 122.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 271.586 123.15 272.734 ;
      VIA 122.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 261.506 123.15 262.654 ;
      VIA 122.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 9.506 123.15 10.654 ;
      VIA 122.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 604.226 78.35 605.374 ;
      VIA 77.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 594.146 78.35 595.294 ;
      VIA 77.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 342.146 78.35 343.294 ;
      VIA 77.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 332.066 78.35 333.214 ;
      VIA 77.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 321.986 78.35 323.134 ;
      VIA 77.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 311.906 78.35 313.054 ;
      VIA 77.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 301.826 78.35 302.974 ;
      VIA 77.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 291.746 78.35 292.894 ;
      VIA 77.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 281.666 78.35 282.814 ;
      VIA 77.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 271.586 78.35 272.734 ;
      VIA 77.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 261.506 78.35 262.654 ;
      VIA 77.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 9.506 78.35 10.654 ;
      VIA 77.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 604.226 33.55 605.374 ;
      VIA 32.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 594.146 33.55 595.294 ;
      VIA 32.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 342.146 33.55 343.294 ;
      VIA 32.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 332.066 33.55 333.214 ;
      VIA 32.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 321.986 33.55 323.134 ;
      VIA 32.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 311.906 33.55 313.054 ;
      VIA 32.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 301.826 33.55 302.974 ;
      VIA 32.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 291.746 33.55 292.894 ;
      VIA 32.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 281.666 33.55 282.814 ;
      VIA 32.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 271.586 33.55 272.734 ;
      VIA 32.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 261.506 33.55 262.654 ;
      VIA 32.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 9.506 33.55 10.654 ;
      VIA 32.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 15.556 595.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 595.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 595.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 595.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 595.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 594.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 594.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 594.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 594.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 594.336 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 594.146 16.19 595.294 ;
      VIA 15.376 595.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 595.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 595.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 595.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 595.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 594.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 594.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 594.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 594.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 594.72 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 585.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 585.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 585.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 585.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 585.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 584.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 584.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 584.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 584.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 584.256 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 584.066 16.19 585.214 ;
      VIA 15.376 585.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 585.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 585.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 585.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 585.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 584.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 584.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 584.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 584.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 584.64 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 574.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 574.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 574.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 574.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 574.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 574.176 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 573.986 16.19 575.134 ;
      VIA 15.376 574.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 574.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 574.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 574.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 574.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 574.56 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 564.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 564.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 564.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 564.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 564.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 564.096 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 563.906 16.19 565.054 ;
      VIA 15.376 564.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 564.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 564.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 564.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 564.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 564.48 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 554.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 554.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 554.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 554.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 554.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 554.016 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 553.826 16.19 554.974 ;
      VIA 15.376 554.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 554.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 554.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 554.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 554.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 554.4 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 544.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 544.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 544.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 544.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 544.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 544.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 544.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 544.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 544.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 544.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 543.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 543.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 543.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 543.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 543.936 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 543.746 16.19 544.894 ;
      VIA 15.376 544.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 544.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 544.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 544.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 544.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 544.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 544.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 544.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 544.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 543.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 543.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 543.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 543.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 543.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 544.32 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 534.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 534.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 534.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 534.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 534.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 534.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 534.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 534.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 534.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 534.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 534.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 534.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 534.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 534.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 534.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 534.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 534.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 534.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 534.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 534.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 534.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 534.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 534.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 534.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 534.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 533.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 533.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 533.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 533.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 533.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 533.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 533.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 533.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 533.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 533.856 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 533.666 16.19 534.814 ;
      VIA 15.376 534.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 534.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 534.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 534.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 534.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 534.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 534.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 534.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 534.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 534.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 534.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 534.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 534.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 534.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 534.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 534.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 534.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 534.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 534.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 534.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 533.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 533.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 533.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 533.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 533.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 533.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 533.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 533.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 533.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 533.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 534.24 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 524.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 524.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 524.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 524.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 524.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 524.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 524.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 524.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 524.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 524.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 524.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 524.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 524.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 524.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 524.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 524.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 524.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 524.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 524.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 524.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 524.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 524.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 524.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 524.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 524.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 523.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 523.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 523.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 523.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 523.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 523.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 523.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 523.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 523.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 523.776 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 523.586 16.19 524.734 ;
      VIA 15.376 524.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 524.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 524.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 524.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 524.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 524.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 524.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 524.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 524.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 524.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 524.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 524.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 524.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 524.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 524.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 524.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 524.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 524.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 524.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 524.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 523.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 523.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 523.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 523.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 523.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 523.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 523.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 523.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 523.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 523.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 524.16 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 514.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 514.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 514.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 514.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 514.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 514.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 514.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 514.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 514.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 514.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 514.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 514.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 514.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 514.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 514.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 514.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 514.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 514.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 514.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 514.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 513.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 513.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 513.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 513.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 513.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 513.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 513.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 513.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 513.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 513.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 513.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 513.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 513.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 513.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 513.696 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 513.506 16.19 514.654 ;
      VIA 15.376 514.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 514.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 514.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 514.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 514.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 514.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 514.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 514.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 514.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 514.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 514.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 514.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 514.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 514.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 514.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 514.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 514.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 514.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 514.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 514.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 513.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 513.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 513.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 513.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 513.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 513.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 513.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 513.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 513.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 513.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 513.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 513.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 513.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 513.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 513.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 514.08 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 504.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 504.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 504.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 504.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 504.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 504.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 504.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 504.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 504.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 504.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 504.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 504.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 504.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 504.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 504.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 503.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 503.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 503.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 503.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 503.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 503.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 503.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 503.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 503.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 503.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 503.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 503.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 503.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 503.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 503.616 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 503.426 16.19 504.574 ;
      VIA 15.376 504.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 504.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 504.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 504.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 504.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 504.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 504.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 504.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 504.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 504.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 504.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 504.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 504.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 504.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 504.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 503.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 503.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 503.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 503.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 503.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 503.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 503.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 503.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 503.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 503.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 503.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 503.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 503.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 503.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 503.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 504 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 494.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 494.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 494.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 494.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 494.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 494.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 494.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 494.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 494.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 494.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 494.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 494.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 494.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 494.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 494.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 493.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 493.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 493.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 493.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 493.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 493.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 493.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 493.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 493.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 493.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 493.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 493.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 493.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 493.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 493.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 493.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 493.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 493.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 493.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 493.536 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 493.346 16.19 494.494 ;
      VIA 15.376 494.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 494.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 494.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 494.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 494.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 494.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 494.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 494.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 494.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 494.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 494.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 494.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 494.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 494.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 494.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 493.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 493.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 493.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 493.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 493.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 493.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 493.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 493.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 493.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 493.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 493.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 493.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 493.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 493.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 493.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 493.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 493.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 493.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 493.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 493.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 493.92 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 484.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 484.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 484.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 484.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 484.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 484.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 484.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 484.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 484.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 484.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 483.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 483.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 483.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 483.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 483.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 483.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 483.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 483.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 483.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 483.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 483.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 483.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 483.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 483.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 483.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 483.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 483.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 483.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 483.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 483.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 483.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 483.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 483.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 483.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 483.456 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 483.266 16.19 484.414 ;
      VIA 15.376 484.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 484.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 484.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 484.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 484.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 484.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 484.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 484.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 484.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 484.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 483.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 483.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 483.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 483.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 483.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 483.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 483.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 483.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 483.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 483.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 483.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 483.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 483.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 483.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 483.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 483.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 483.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 483.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 483.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 483.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 483.84 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 474.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 474.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 474.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 474.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 474.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 474.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 474.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 474.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 474.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 474.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 473.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 473.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 473.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 473.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 473.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 473.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 473.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 473.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 473.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 473.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 473.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 473.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 473.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 473.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 473.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 473.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 473.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 473.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 473.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 473.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 473.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 473.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 473.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 473.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 473.376 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 473.186 16.19 474.334 ;
      VIA 15.376 474.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 474.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 474.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 474.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 474.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 474.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 474.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 474.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 474.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 474.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 473.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 473.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 473.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 473.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 473.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 473.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 473.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 473.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 473.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 473.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 473.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 473.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 473.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 473.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 473.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 473.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 473.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 473.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 473.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 473.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 473.76 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 464.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 464.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 464.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 464.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 464.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 463.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 463.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 463.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 463.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 463.296 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 463.106 16.19 464.254 ;
      VIA 15.376 464.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 464.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 464.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 464.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 464.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 463.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 463.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 463.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 463.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 463.68 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 453.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 453.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 453.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 453.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 453.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 453.216 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 453.026 16.19 454.174 ;
      VIA 15.376 453.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 453.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 453.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 453.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 453.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 453.6 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 443.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 443.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 443.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 443.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 443.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 443.136 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 442.946 16.19 444.094 ;
      VIA 15.376 443.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 443.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 443.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 443.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 443.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 443.52 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 433.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 433.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 433.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 433.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 433.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 433.056 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 432.866 16.19 434.014 ;
      VIA 15.376 433.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 433.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 433.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 433.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 433.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 433.44 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 423.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 423.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 423.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 423.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 423.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 423.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 423.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 423.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 423.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 423.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 422.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 422.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 422.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 422.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 422.976 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 422.786 16.19 423.934 ;
      VIA 15.376 423.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 423.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 423.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 423.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 423.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 423.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 423.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 423.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 423.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 422.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 422.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 422.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 422.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 422.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 423.36 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 413.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 413.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 413.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 413.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 413.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 413.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 413.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 413.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 413.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 413.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 412.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 412.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 412.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 412.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 412.896 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 412.706 16.19 413.854 ;
      VIA 15.376 413.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 413.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 413.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 413.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 413.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 413.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 413.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 413.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 413.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 412.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 412.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 412.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 412.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 412.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 413.28 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 403.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 403.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 403.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 403.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 403.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 403.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 403.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 403.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 403.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 403.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 403.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 403.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 403.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 403.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 403.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 403.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 403.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 403.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 403.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 403.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 403.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 403.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 403.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 403.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 403.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 402.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 402.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 402.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 402.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 402.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 402.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 402.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 402.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 402.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 402.816 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 402.626 16.19 403.774 ;
      VIA 15.376 403.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 403.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 403.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 403.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 403.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 403.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 403.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 403.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 403.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 403.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 403.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 403.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 403.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 403.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 403.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 403.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 403.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 403.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 403.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 403.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 402.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 402.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 402.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 402.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 402.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 402.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 402.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 402.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 402.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 402.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 403.2 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 393.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 393.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 393.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 393.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 393.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 393.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 393.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 393.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 393.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 393.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 393.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 393.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 393.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 393.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 393.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 393.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 393.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 393.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 393.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 393.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 392.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 392.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 392.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 392.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 392.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 392.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 392.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 392.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 392.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 392.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 392.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 392.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 392.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 392.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 392.736 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 392.546 16.19 393.694 ;
      VIA 15.376 393.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 393.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 393.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 393.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 393.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 393.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 393.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 393.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 393.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 393.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 393.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 393.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 393.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 393.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 393.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 393.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 393.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 393.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 393.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 393.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 392.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 392.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 392.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 392.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 392.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 392.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 392.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 392.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 392.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 392.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 392.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 392.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 392.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 392.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 392.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 393.12 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 383.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 383.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 383.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 383.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 383.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 383.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 383.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 383.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 383.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 383.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 383.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 383.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 383.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 383.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 383.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 383.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 383.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 383.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 383.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 383.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 382.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 382.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 382.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 382.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 382.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 382.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 382.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 382.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 382.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 382.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 382.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 382.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 382.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 382.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 382.656 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 382.466 16.19 383.614 ;
      VIA 15.376 383.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 383.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 383.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 383.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 383.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 383.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 383.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 383.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 383.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 383.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 383.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 383.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 383.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 383.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 383.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 383.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 383.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 383.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 383.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 383.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 382.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 382.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 382.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 382.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 382.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 382.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 382.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 382.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 382.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 382.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 382.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 382.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 382.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 382.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 382.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 383.04 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 373.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 373.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 373.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 373.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 373.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 373.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 373.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 373.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 373.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 373.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 373.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 373.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 373.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 373.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 373.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 372.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 372.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 372.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 372.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 372.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 372.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 372.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 372.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 372.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 372.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 372.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 372.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 372.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 372.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 372.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 372.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 372.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 372.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 372.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 372.576 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 372.386 16.19 373.534 ;
      VIA 15.376 373.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 373.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 373.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 373.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 373.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 373.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 373.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 373.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 373.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 373.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 373.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 373.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 373.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 373.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 373.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 372.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 372.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 372.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 372.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 372.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 372.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 372.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 372.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 372.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 372.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 372.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 372.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 372.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 372.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 372.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 372.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 372.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 372.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 372.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 372.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 372.96 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 363.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 363.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 363.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 363.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 363.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 363.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 363.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 363.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 363.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 363.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 363.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 363.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 363.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 363.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 363.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 362.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 362.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 362.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 362.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 362.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 362.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 362.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 362.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 362.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 362.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 362.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 362.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 362.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 362.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 362.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 362.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 362.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 362.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 362.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 362.496 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 362.306 16.19 363.454 ;
      VIA 15.376 363.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 363.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 363.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 363.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 363.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 363.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 363.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 363.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 363.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 363.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 363.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 363.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 363.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 363.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 363.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 362.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 362.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 362.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 362.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 362.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 362.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 362.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 362.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 362.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 362.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 362.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 362.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 362.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 362.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 362.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 362.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 362.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 362.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 362.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 362.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 362.88 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 353.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 353.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 353.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 353.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 353.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 353.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 353.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 353.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 353.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 353.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 352.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 352.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 352.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 352.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 352.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 352.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 352.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 352.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 352.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 352.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 352.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 352.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 352.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 352.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 352.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 352.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 352.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 352.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 352.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 352.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 352.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 352.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 352.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 352.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 352.416 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 352.226 16.19 353.374 ;
      VIA 15.376 353.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 353.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 353.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 353.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 353.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 353.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 353.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 353.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 353.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 353.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 352.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 352.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 352.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 352.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 352.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 352.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 352.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 352.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 352.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 352.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 352.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 352.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 352.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 352.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 352.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 352.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 352.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 352.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 352.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 352.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 352.8 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 343.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 343.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 343.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 343.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 343.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 342.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 342.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 342.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 342.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 342.336 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 342.146 16.19 343.294 ;
      VIA 15.376 343.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 343.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 343.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 343.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 343.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 342.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 342.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 342.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 342.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 342.72 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 262.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 262.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 262.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 262.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 262.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 262.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 262.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 262.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 262.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 262.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 262.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 262.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 262.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 262.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 262.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 262.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 262.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 262.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 262.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 262.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 261.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 261.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 261.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 261.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 261.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 261.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 261.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 261.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 261.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 261.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 261.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 261.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 261.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 261.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 261.696 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 261.506 16.19 262.654 ;
      VIA 15.376 262.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 262.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 262.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 262.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 262.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 262.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 262.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 262.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 262.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 262.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 262.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 262.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 262.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 262.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 262.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 262.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 262.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 262.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 262.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 262.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 261.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 261.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 261.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 261.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 261.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 261.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 261.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 261.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 261.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 261.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 261.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 261.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 261.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 261.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 261.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 262.08 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 252.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 252.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 252.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 252.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 252.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 252.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 252.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 252.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 252.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 252.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 252.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 252.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 252.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 252.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 252.128 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 252 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 252 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 252 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 252 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 252 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 251.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 251.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 251.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 251.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 251.872 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 251.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 251.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 251.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 251.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 251.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 251.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 251.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 251.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 251.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 251.616 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 251.426 16.19 252.574 ;
      VIA 15.376 252.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 252.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 252.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 252.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 252.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 252.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 252.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 252.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 252.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 252.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 252.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 252.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 252.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 252.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 252.128 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 252 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 252 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 252 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 252 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 252 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 251.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 251.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 251.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 251.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 251.872 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 251.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 251.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 251.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 251.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 251.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 251.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 251.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 251.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 251.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 251.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 252 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 242.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 242.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 242.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 242.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 242.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 242.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 242.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 242.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 242.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 242.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 242.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 242.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 242.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 242.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 242.048 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 241.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 241.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 241.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 241.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 241.92 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 241.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 241.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 241.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 241.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 241.792 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 241.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 241.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 241.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 241.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 241.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 241.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 241.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 241.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 241.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 241.536 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 241.346 16.19 242.494 ;
      VIA 15.376 242.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 242.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 242.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 242.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 242.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 242.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 242.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 242.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 242.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 242.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 242.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 242.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 242.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 242.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 242.048 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 241.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 241.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 241.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 241.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 241.92 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 241.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 241.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 241.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 241.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 241.792 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 241.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 241.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 241.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 241.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 241.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 241.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 241.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 241.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 241.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 241.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 241.92 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 232.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 232.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 232.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 232.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 232.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 232.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 232.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 232.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 232.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 232.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 231.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 231.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 231.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 231.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 231.968 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 231.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 231.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 231.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 231.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 231.84 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 231.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 231.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 231.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 231.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 231.712 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 231.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 231.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 231.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 231.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 231.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 231.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 231.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 231.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 231.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 231.456 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 231.266 16.19 232.414 ;
      VIA 15.376 232.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 232.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 232.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 232.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 232.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 232.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 232.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 232.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 232.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 232.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 231.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 231.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 231.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 231.968 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 231.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 231.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 231.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 231.84 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 231.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 231.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 231.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 231.712 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 231.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 231.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 231.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 231.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 231.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 231.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 231.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 231.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 231.84 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 222.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 222.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 222.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 222.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 222.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 222.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 222.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 222.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 222.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 222.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 221.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 221.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 221.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 221.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 221.888 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 221.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 221.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 221.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 221.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 221.76 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 221.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 221.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 221.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 221.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 221.632 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 221.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 221.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 221.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 221.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 221.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 221.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 221.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 221.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 221.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 221.376 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 221.186 16.19 222.334 ;
      VIA 15.376 222.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 222.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 222.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 222.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 222.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 222.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 222.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 222.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 222.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 222.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 221.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 221.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 221.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 221.888 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 221.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 221.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 221.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 221.76 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 221.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 221.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 221.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 221.632 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 221.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 221.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 221.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 221.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 221.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 221.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 221.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 221.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 221.76 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 212.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 212.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 212.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 212.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 212.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.808 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.68 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.552 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 211.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 211.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 211.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 211.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 211.296 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 211.106 16.19 212.254 ;
      VIA 15.376 212.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 212.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 212.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 212.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 212.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.808 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.68 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.552 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 211.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 211.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 211.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 211.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 211.68 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 201.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.728 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.6 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.472 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 201.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 201.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 201.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 201.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 201.216 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 201.026 16.19 202.174 ;
      VIA 15.376 201.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.728 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.6 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.472 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 201.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 201.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 201.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 201.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 201.6 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 191.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.648 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.52 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.392 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 191.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 191.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 191.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 191.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 191.136 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 190.946 16.19 192.094 ;
      VIA 15.376 191.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.648 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.52 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.392 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 191.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 191.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 191.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 191.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 191.52 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 181.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.568 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.44 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.312 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 181.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 181.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 181.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 181.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 181.056 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 180.866 16.19 182.014 ;
      VIA 15.376 181.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.568 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.44 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.312 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 181.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 181.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 181.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 181.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 181.44 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 171.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.744 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 171.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.616 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 171.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.488 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 171.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.36 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 171.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.232 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 171.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 171.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 171.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 171.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 171.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 170.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 170.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 170.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 170.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 170.976 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 170.786 16.19 171.934 ;
      VIA 15.376 171.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.744 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 171.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.616 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 171.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.488 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 171.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.36 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 171.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.232 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 171.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 171.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 171.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 171.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 170.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 170.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 170.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 170.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 170.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 171.36 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 161.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.664 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 161.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.536 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 161.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.408 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 161.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.28 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 161.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.152 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 161.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 161.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 161.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 161.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 161.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 160.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 160.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 160.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 160.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 160.896 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 160.706 16.19 161.854 ;
      VIA 15.376 161.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.664 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 161.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.536 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 161.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.408 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 161.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.28 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 161.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.152 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 161.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 161.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 161.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 161.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 160.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 160.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 160.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 160.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 160.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 161.28 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 151.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 151.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 151.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 151.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 151.584 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 151.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 151.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 151.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 151.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 151.456 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 151.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 151.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 151.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 151.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 151.328 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 151.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 151.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 151.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 151.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 151.2 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 151.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 151.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 151.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 151.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 151.072 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 150.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 150.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 150.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 150.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 150.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 150.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 150.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 150.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 150.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 150.816 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 150.626 16.19 151.774 ;
      VIA 15.376 151.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 151.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 151.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 151.584 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 151.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 151.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 151.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 151.456 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 151.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 151.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 151.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 151.328 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 151.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 151.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 151.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 151.2 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 151.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 151.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 151.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 151.072 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 150.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 150.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 150.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 150.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 150.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 150.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 150.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 150.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 150.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 150.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 151.2 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 141.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 141.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 141.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 141.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 141.504 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 141.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 141.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 141.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 141.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 141.376 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 141.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 141.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 141.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 141.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 141.248 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 141.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 141.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 141.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 141.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 141.12 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 140.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 140.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 140.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 140.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 140.992 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 140.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 140.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 140.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 140.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 140.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 140.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 140.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 140.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 140.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 140.736 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 140.546 16.19 141.694 ;
      VIA 15.376 141.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 141.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 141.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 141.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 141.504 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 141.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 141.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 141.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 141.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 141.376 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 141.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 141.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 141.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 141.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 141.248 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 141.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 141.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 141.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 141.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 141.12 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 140.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 140.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 140.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 140.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 140.992 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 140.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 140.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 140.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 140.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 140.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 140.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 140.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 140.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 140.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 140.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 141.12 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 131.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 131.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 131.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 131.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 131.424 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 131.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 131.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 131.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 131.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 131.296 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 131.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 131.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 131.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 131.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 131.168 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 131.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 131.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 131.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 131.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 131.04 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 130.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 130.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 130.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 130.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 130.912 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 130.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 130.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 130.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 130.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 130.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 130.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 130.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 130.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 130.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 130.656 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 130.466 16.19 131.614 ;
      VIA 15.376 131.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 131.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 131.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 131.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 131.424 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 131.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 131.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 131.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 131.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 131.296 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 131.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 131.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 131.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 131.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 131.168 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 131.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 131.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 131.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 131.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 131.04 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 130.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 130.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 130.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 130.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 130.912 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 130.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 130.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 130.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 130.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 130.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 130.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 130.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 130.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 130.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 130.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 131.04 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 121.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 121.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 121.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 121.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 121.344 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 121.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 121.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 121.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 121.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 121.216 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 121.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 121.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 121.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 121.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 121.088 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 120.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 120.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 120.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 120.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 120.96 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 120.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 120.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 120.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 120.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 120.832 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 120.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 120.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 120.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 120.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 120.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 120.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 120.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 120.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 120.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 120.576 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 120.386 16.19 121.534 ;
      VIA 15.376 121.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 121.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 121.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 121.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 121.344 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 121.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 121.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 121.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 121.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 121.216 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 121.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 121.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 121.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 121.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 121.088 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 120.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 120.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 120.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 120.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 120.96 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 120.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 120.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 120.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 120.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 120.832 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 120.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 120.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 120.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 120.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 120.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 120.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 120.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 120.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 120.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 120.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 120.96 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 111.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 111.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 111.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 111.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 111.264 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 111.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 111.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 111.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 111.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 111.136 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 111.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 111.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 111.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 111.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 111.008 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 110.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 110.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 110.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 110.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 110.88 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 110.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 110.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 110.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 110.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 110.752 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 110.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 110.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 110.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 110.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 110.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 110.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 110.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 110.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 110.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 110.496 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 110.306 16.19 111.454 ;
      VIA 15.376 111.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 111.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 111.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 111.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 111.264 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 111.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 111.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 111.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 111.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 111.136 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 111.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 111.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 111.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 111.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 111.008 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 110.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 110.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 110.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 110.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 110.88 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 110.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 110.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 110.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 110.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 110.752 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 110.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 110.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 110.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 110.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 110.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 110.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 110.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 110.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 110.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 110.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 110.88 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 101.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 101.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 101.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 101.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 101.184 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 101.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 101.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 101.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 101.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 101.056 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 100.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 100.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 100.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 100.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 100.928 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 100.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 100.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 100.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 100.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 100.8 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 100.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 100.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 100.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 100.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 100.672 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 100.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 100.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 100.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 100.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 100.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 100.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 100.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 100.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 100.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 100.416 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 100.226 16.19 101.374 ;
      VIA 15.376 101.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 101.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 101.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 101.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 101.184 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 101.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 101.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 101.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 101.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 101.056 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 100.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 100.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 100.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 100.928 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 100.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 100.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 100.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 100.8 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 100.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 100.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 100.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 100.672 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 100.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 100.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 100.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 100.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 100.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 100.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 100.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 100.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 100.8 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 91.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 91.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 91.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 91.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 91.104 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.976 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.848 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.72 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.592 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 90.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 90.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 90.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 90.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 90.336 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 90.146 16.19 91.294 ;
      VIA 15.376 91.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 91.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 91.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 91.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 91.104 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.976 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.848 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.72 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.592 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 90.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 90.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 90.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 90.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 90.72 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 81.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 81.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 81.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 81.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 81.024 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.896 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.768 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.64 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.512 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.384 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 80.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 80.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 80.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 80.256 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 80.256 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 80.066 16.19 81.214 ;
      VIA 15.376 81.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 81.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 81.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 81.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 81.024 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.896 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.768 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.64 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.512 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.384 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 80.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 80.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 80.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 80.256 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 80.64 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 70.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.944 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.816 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.688 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.56 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.432 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.304 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 70.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 70.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 70.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 70.176 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 70.176 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 69.986 16.19 71.134 ;
      VIA 15.376 70.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.944 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.816 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.688 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.56 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.432 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.304 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 70.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 70.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 70.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 70.176 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 70.56 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 60.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.864 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.736 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.608 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.48 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.352 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.224 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 60.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 60.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 60.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 60.096 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 60.096 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 59.906 16.19 61.054 ;
      VIA 15.376 60.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.864 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.736 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.608 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.48 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.352 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.224 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 60.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 60.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 60.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 60.096 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 60.48 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 50.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.784 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.656 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.528 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.4 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.272 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.144 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 50.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 50.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 50.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 50.016 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 50.016 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 49.826 16.19 50.974 ;
      VIA 15.376 50.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.784 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.656 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.528 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.4 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.272 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.144 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 50.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 50.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 50.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 50.016 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 50.4 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 40.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.704 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 40.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.576 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 40.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.448 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 40.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.32 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 40.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.192 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 40.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 40.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 40.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 40.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 40.064 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 39.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 39.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 39.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 39.936 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 39.936 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 39.746 16.19 40.894 ;
      VIA 15.376 40.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.704 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 40.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.576 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 40.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.448 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 40.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.32 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 40.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.192 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 40.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 40.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 40.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 40.064 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 39.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 39.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 39.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 39.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 39.936 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 40.32 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 30.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 30.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 30.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 30.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 30.624 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 30.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 30.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 30.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 30.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 30.496 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 30.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 30.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 30.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 30.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 30.368 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 30.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 30.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 30.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 30.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 30.24 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 30.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 30.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 30.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 30.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 30.112 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 29.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 29.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 29.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 29.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 29.984 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 29.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 29.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 29.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 29.856 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 29.856 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 29.666 16.19 30.814 ;
      VIA 15.376 30.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 30.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 30.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 30.624 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 30.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 30.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 30.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 30.496 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 30.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 30.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 30.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 30.368 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 30.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 30.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 30.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 30.24 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 30.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 30.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 30.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 30.112 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 29.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 29.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 29.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 29.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 29.984 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 29.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 29.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 29.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 29.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 29.856 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 30.24 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 20.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 20.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 20.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 20.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 20.544 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 20.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 20.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 20.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 20.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 20.416 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 20.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 20.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 20.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 20.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 20.288 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 20.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 20.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 20.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 20.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 20.16 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 20.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 20.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 20.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 20.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 20.032 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 19.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 19.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 19.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 19.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 19.904 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 19.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 19.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 19.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 19.776 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 19.776 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 19.586 16.19 20.734 ;
      VIA 15.376 20.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 20.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 20.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 20.544 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 20.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 20.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 20.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 20.416 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 20.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 20.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 20.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 20.288 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 20.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 20.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 20.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 20.16 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 20.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 20.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 20.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 20.032 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 19.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 19.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 19.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 19.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 19.904 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 19.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 19.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 19.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 19.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 19.776 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 20.16 via1_2_4480_1800_1_4_1240_1240 ;
      VIA 15.556 10.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 10.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 10.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 10.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 10.464 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 10.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 10.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 10.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 10.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 10.336 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 10.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 10.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 10.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 10.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 10.208 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 10.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 10.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 10.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 10.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 10.08 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 9.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 9.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 9.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 9.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 9.952 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 9.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 9.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 9.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 9.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 9.824 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.556 9.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.428 9.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.3 9.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.172 9.696 via3_4_4480_1800_1_1_256_256 ;
      VIA 15.044 9.696 via3_4_4480_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  14.05 9.506 16.19 10.654 ;
      VIA 15.376 10.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 10.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 10.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 10.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 10.464 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 10.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 10.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 10.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 10.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 10.336 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 10.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 10.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 10.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 10.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 10.208 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 10.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 10.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 10.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 10.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 10.08 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 9.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 9.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 9.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 9.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 9.952 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 9.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 9.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 9.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 9.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 9.824 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.376 9.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.248 9.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 9.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.992 9.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 14.864 9.696 via2_3_4480_1800_1_1_256_256 ;
      VIA 15.12 10.08 via1_2_4480_1800_1_4_1240_1240 ;
    END
  END VSS
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  360.68 0 361.12 1.28 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  362.48 0 362.92 1.28 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  175.28 0 175.72 1.28 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  364.28 0 364.72 1.28 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  366.08 0 366.52 1.28 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  367.88 0 368.32 1.28 ;
    END
  END addr[5]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  369.68 0 370.12 1.28 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  160.88 0 161.32 1.28 ;
    END
  END clk
  PIN idat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 19.46 0.52 19.74 ;
    END
  END idat[0]
  PIN idat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 357.7 0.52 357.98 ;
    END
  END idat[10]
  PIN idat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 347.62 0.52 347.9 ;
    END
  END idat[11]
  PIN idat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 353.22 0.52 353.5 ;
    END
  END idat[12]
  PIN idat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  378.68 618.72 379.12 620 ;
    END
  END idat[13]
  PIN idat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  385.88 618.72 386.32 620 ;
    END
  END idat[14]
  PIN idat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  438.08 618.72 438.52 620 ;
    END
  END idat[15]
  PIN idat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  560.48 0 560.92 1.28 ;
    END
  END idat[16]
  PIN idat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  612.68 0 613.12 1.28 ;
    END
  END idat[17]
  PIN idat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  618.08 0 618.52 1.28 ;
    END
  END idat[18]
  PIN idat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  670.28 0 670.72 1.28 ;
    END
  END idat[19]
  PIN idat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  81.68 0 82.12 1.28 ;
    END
  END idat[1]
  PIN idat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  859.28 0 859.72 1.28 ;
    END
  END idat[20]
  PIN idat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  909.68 0 910.12 1.28 ;
    END
  END idat[21]
  PIN idat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  916.88 0 917.32 1.28 ;
    END
  END idat[22]
  PIN idat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  969.08 0 969.52 1.28 ;
    END
  END idat[23]
  PIN idat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  560.48 618.72 560.92 620 ;
    END
  END idat[24]
  PIN idat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  612.68 618.72 613.12 620 ;
    END
  END idat[25]
  PIN idat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  618.08 618.72 618.52 620 ;
    END
  END idat[26]
  PIN idat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 357.7 1020 357.98 ;
    END
  END idat[27]
  PIN idat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 356.58 1020 356.86 ;
    END
  END idat[28]
  PIN idat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 355.46 1020 355.74 ;
    END
  END idat[29]
  PIN idat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  87.08 0 87.52 1.28 ;
    END
  END idat[2]
  PIN idat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 353.22 1020 353.5 ;
    END
  END idat[30]
  PIN idat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 349.86 1020 350.14 ;
    END
  END idat[31]
  PIN idat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  139.28 0 139.72 1.28 ;
    END
  END idat[3]
  PIN idat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  328.28 0 328.72 1.28 ;
    END
  END idat[4]
  PIN idat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  378.68 0 379.12 1.28 ;
    END
  END idat[5]
  PIN idat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  385.88 0 386.32 1.28 ;
    END
  END idat[6]
  PIN idat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  438.08 0 438.52 1.28 ;
    END
  END idat[7]
  PIN idat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 350.98 0.52 351.26 ;
    END
  END idat[8]
  PIN idat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 355.46 0.52 355.74 ;
    END
  END idat[9]
  PIN odat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 20.58 0.52 20.86 ;
    END
  END odat[0]
  PIN odat[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 348.74 0.52 349.02 ;
    END
  END odat[10]
  PIN odat[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 352.1 0.52 352.38 ;
    END
  END odat[11]
  PIN odat[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 354.34 0.52 354.62 ;
    END
  END odat[12]
  PIN odat[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  375.08 618.72 375.52 620 ;
    END
  END odat[13]
  PIN odat[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  389.48 618.72 389.92 620 ;
    END
  END odat[14]
  PIN odat[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  429.08 618.72 429.52 620 ;
    END
  END odat[15]
  PIN odat[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  567.68 0 568.12 1.28 ;
    END
  END odat[16]
  PIN odat[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  609.08 0 609.52 1.28 ;
    END
  END odat[17]
  PIN odat[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  621.68 0 622.12 1.28 ;
    END
  END odat[18]
  PIN odat[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  663.08 0 663.52 1.28 ;
    END
  END odat[19]
  PIN odat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  78.08 0 78.52 1.28 ;
    END
  END odat[1]
  PIN odat[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  866.48 0 866.92 1.28 ;
    END
  END odat[20]
  PIN odat[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  906.08 0 906.52 1.28 ;
    END
  END odat[21]
  PIN odat[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  920.48 0 920.92 1.28 ;
    END
  END odat[22]
  PIN odat[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  960.08 0 960.52 1.28 ;
    END
  END odat[23]
  PIN odat[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  567.68 618.72 568.12 620 ;
    END
  END odat[24]
  PIN odat[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  609.08 618.72 609.52 620 ;
    END
  END odat[25]
  PIN odat[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  621.68 618.72 622.12 620 ;
    END
  END odat[26]
  PIN odat[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 352.1 1020 352.38 ;
    END
  END odat[27]
  PIN odat[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 350.98 1020 351.26 ;
    END
  END odat[28]
  PIN odat[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 354.34 1020 354.62 ;
    END
  END odat[29]
  PIN odat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  90.68 0 91.12 1.28 ;
    END
  END odat[2]
  PIN odat[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 348.74 1020 349.02 ;
    END
  END odat[30]
  PIN odat[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  1019.48 347.62 1020 347.9 ;
    END
  END odat[31]
  PIN odat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  132.08 0 132.52 1.28 ;
    END
  END odat[3]
  PIN odat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  335.48 0 335.92 1.28 ;
    END
  END odat[4]
  PIN odat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  375.08 0 375.52 1.28 ;
    END
  END odat[5]
  PIN odat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  389.48 0 389.92 1.28 ;
    END
  END odat[6]
  PIN odat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  429.08 0 429.52 1.28 ;
    END
  END odat[7]
  PIN odat[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 356.58 0.52 356.86 ;
    END
  END odat[8]
  PIN odat[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 349.86 0.52 350.14 ;
    END
  END odat[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  488.48 0 488.92 1.28 ;
    END
  END we
  OBS
    LAYER Metal1 ;
     RECT  10.08 9.63 13.325 610.29 ;
     RECT  13.325 8.845 16.685 610.29 ;
     RECT  16.685 7.725 160.275 610.29 ;
     RECT  160.275 8.285 191.635 610.29 ;
     RECT  191.635 9.63 272.045 610.29 ;
     RECT  272.045 6.605 296.685 610.29 ;
     RECT  296.685 6.045 416.755 610.29 ;
     RECT  416.755 6.605 453.715 610.29 ;
     RECT  453.715 7.165 541.965 610.29 ;
     RECT  541.965 6.605 544.205 610.29 ;
     RECT  544.205 5.485 706.275 610.29 ;
     RECT  706.275 6.045 714.115 610.29 ;
     RECT  714.115 6.605 722.515 610.29 ;
     RECT  722.515 7.165 803.155 610.29 ;
     RECT  803.155 9.63 906.525 610.29 ;
     RECT  906.525 8.845 944.835 610.29 ;
     RECT  944.835 9.63 960.285 610.29 ;
     RECT  960.285 8.285 966.115 610.29 ;
     RECT  966.115 9.63 1009.68 610.29 ;
    LAYER Metal2 ;
     RECT  544.18 5.46 544.46 6.02 ;
     RECT  706.02 5.46 706.3 6.02 ;
     RECT  544.18 6.02 546.14 6.58 ;
     RECT  706.02 6.02 714.14 6.58 ;
     RECT  296.66 6.02 296.94 7.14 ;
     RECT  358.26 6.58 358.54 7.14 ;
     RECT  541.94 6.58 546.14 7.14 ;
     RECT  380.1 7.14 380.38 7.7 ;
     RECT  462.98 7.14 463.26 7.7 ;
     RECT  541.94 7.14 550.62 7.7 ;
     RECT  613.06 7.7 623.98 8.07 ;
     RECT  16.66 7.7 16.94 8.26 ;
     RECT  68.74 7.14 69.02 8.26 ;
     RECT  347.62 7.14 358.54 8.26 ;
     RECT  380.1 7.7 383.74 8.26 ;
     RECT  404.74 7.14 405.02 8.26 ;
     RECT  571.06 8.07 571.34 8.26 ;
     RECT  663.46 8.07 663.74 8.26 ;
     RECT  960.26 8.07 960.54 8.26 ;
     RECT  176.26 8.26 176.54 8.63 ;
     RECT  191.38 8.26 191.66 8.63 ;
     RECT  16.66 8.26 19.74 8.82 ;
     RECT  292.74 7.14 296.94 8.82 ;
     RECT  462.98 7.7 463.82 8.82 ;
     RECT  609.14 8.07 623.98 8.82 ;
     RECT  906.5 8.63 906.78 8.82 ;
     RECT  923.86 8.63 924.14 8.82 ;
     RECT  68.74 8.26 72.94 9.38 ;
     RECT  330.82 8.82 332.22 9.38 ;
     RECT  433.3 6.58 434.14 9.38 ;
     RECT  448.98 8.26 449.26 9.38 ;
     RECT  536.34 7.7 550.62 9.38 ;
     RECT  571.06 8.26 576.94 9.38 ;
     RECT  960.26 8.26 966.14 9.38 ;
     RECT  35.7 8.82 39.34 9.506 ;
     RECT  160.02 7.7 160.3 9.506 ;
     RECT  176.26 8.63 191.66 9.506 ;
     RECT  223.3 6.58 223.58 9.506 ;
     RECT  347.62 8.26 405.02 9.506 ;
     RECT  536.34 9.38 576.94 9.506 ;
     RECT  663.46 8.26 669.9 9.506 ;
     RECT  706.02 6.58 722.54 9.506 ;
     RECT  752.5 7.7 752.78 9.506 ;
     RECT  802.9 7.14 803.18 9.506 ;
     RECT  906.5 8.82 924.14 9.506 ;
     RECT  960.26 9.38 970.9 9.506 ;
     RECT  314.865 8.82 315.145 10.5 ;
     RECT  326.62 9.38 332.22 10.5 ;
     RECT  479.41 9.506 481.55 11.025 ;
     RECT  416.5 6.02 416.78 11.06 ;
     RECT  433.3 9.38 449.26 11.06 ;
     RECT  121.01 9.506 123.15 11.34 ;
     RECT  609.14 8.82 629.58 11.34 ;
     RECT  860.3 9.38 860.58 11.34 ;
     RECT  906.5 9.506 929.55 11.34 ;
     RECT  960.26 9.506 974.35 11.34 ;
     RECT  292.74 8.82 303.1 11.62 ;
     RECT  314.865 10.5 332.22 11.62 ;
     RECT  602.765 11.34 629.58 11.62 ;
     RECT  658.61 9.506 669.9 11.62 ;
     RECT  901.805 11.34 929.55 11.62 ;
     RECT  944.58 8.82 944.86 11.62 ;
     RECT  121.01 11.34 128.165 12.18 ;
     RECT  140.14 9.38 140.42 12.18 ;
     RECT  13.02 8.82 19.74 12.31 ;
     RECT  31.41 9.506 39.34 12.31 ;
     RECT  68.74 9.38 82.18 12.31 ;
     RECT  101.445 11.34 105.085 12.31 ;
     RECT  292.74 11.62 332.22 12.31 ;
     RECT  345.01 9.506 405.02 12.31 ;
     RECT  602.765 11.62 630.42 12.31 ;
     RECT  645.54 8.26 645.82 12.31 ;
     RECT  857.565 11.34 860.58 12.31 ;
     RECT  292.74 12.31 405.02 12.46 ;
     RECT  416.5 11.06 449.485 12.46 ;
     RECT  121.01 12.18 140.42 13.02 ;
     RECT  658.61 11.62 673.54 13.02 ;
     RECT  857.565 12.31 870.1 13.02 ;
     RECT  882.61 9.506 884.75 13.02 ;
     RECT  958.365 11.34 974.35 13.02 ;
     RECT  292.74 12.46 449.485 13.3 ;
     RECT  461.86 8.82 463.82 13.3 ;
     RECT  958.365 13.02 976.78 13.3 ;
     RECT  824.18 13.3 825.02 13.86 ;
     RECT  837.81 9.506 839.95 13.86 ;
     RECT  958.365 13.3 983.5 13.86 ;
     RECT  13.02 12.31 39.34 14.546 ;
     RECT  255.41 9.506 257.55 14.546 ;
     RECT  272.02 6.58 272.3 14.546 ;
     RECT  748.21 9.506 752.78 14.546 ;
     RECT  824.18 13.86 839.95 14.546 ;
     RECT  857.565 13.02 884.75 14.546 ;
     RECT  958.365 13.86 984.06 14.546 ;
     RECT  999.09 9.506 1001.23 14.546 ;
     RECT  11.25 14.546 39.34 16.1 ;
     RECT  824.18 14.546 844.99 16.66 ;
     RECT  9.94 16.1 39.34 20 ;
     RECT  62.86 12.31 105.085 20 ;
     RECT  121.01 13.02 146.3 20 ;
     RECT  160.02 9.506 191.66 20 ;
     RECT  210.61 9.506 223.58 20 ;
     RECT  255.41 14.546 272.3 20 ;
     RECT  292.74 13.3 463.82 20 ;
     RECT  524.21 9.506 576.94 20 ;
     RECT  602.765 12.31 645.82 20 ;
     RECT  658.61 13.02 679.42 20 ;
     RECT  690.9 7.7 691.18 20 ;
     RECT  703.41 9.506 722.54 20 ;
     RECT  748.21 14.546 755.39 20 ;
     RECT  793.01 9.506 803.18 20 ;
     RECT  823.9 16.66 844.99 20 ;
     RECT  857.565 14.546 889.79 20 ;
     RECT  901.805 11.62 944.86 20 ;
     RECT  958.365 14.546 1001.23 20 ;
     RECT  479.41 11.025 491.82 41.3 ;
     RECT  479.41 41.3 492.38 59.22 ;
     RECT  479.41 59.22 492.66 62.02 ;
     RECT  479.41 62.02 496.86 62.3 ;
     RECT  479.41 62.3 493.5 63.42 ;
     RECT  9.94 20 463.82 100.94 ;
     RECT  9.94 100.94 462.7 159.46 ;
     RECT  9.94 159.46 463.82 184.1 ;
     RECT  479.41 63.42 486.59 188.58 ;
     RECT  9.94 184.1 466.06 188.86 ;
     RECT  479.41 188.58 490.14 188.86 ;
     RECT  9.94 188.86 486.59 192.78 ;
     RECT  9.94 192.78 465.5 252.88 ;
     RECT  524.21 20 1001.23 252.88 ;
     RECT  972.21 252.88 1001.23 257.614 ;
     RECT  999.09 257.614 1001.23 262.654 ;
     RECT  300.21 252.88 307.39 264.55 ;
     RECT  345.01 252.88 352.19 264.55 ;
     RECT  165.81 252.88 172.99 264.74 ;
     RECT  293.86 264.55 307.39 264.88 ;
     RECT  345.01 264.55 352.94 264.88 ;
     RECT  454.02 252.88 465.5 265.02 ;
     RECT  160.02 264.74 172.99 268.66 ;
     RECT  454.02 265.02 462.7 276.5 ;
     RECT  9.94 252.88 18.62 277.34 ;
     RECT  453.46 276.5 462.7 280.14 ;
     RECT  158.9 268.66 172.99 294.14 ;
     RECT  9.94 277.34 18.06 325.5 ;
     RECT  9.94 325.5 19.045 325.78 ;
     RECT  9.94 325.78 19.18 328.39 ;
     RECT  31.41 252.88 38.59 328.39 ;
     RECT  160.02 294.14 172.99 328.39 ;
     RECT  389.81 252.88 396.99 329.7 ;
     RECT  411.46 329.51 411.74 329.84 ;
     RECT  613.81 252.88 620.99 330.26 ;
     RECT  235.06 328.39 235.34 330.4 ;
     RECT  748.21 252.88 755.39 330.63 ;
     RECT  327.46 329.7 327.74 330.82 ;
     RECT  345.01 264.88 352.19 330.82 ;
     RECT  454.02 280.14 462.7 330.82 ;
     RECT  972.21 257.614 984.62 330.82 ;
     RECT  121.01 252.88 128.19 331.38 ;
     RECT  139.86 330.26 140.14 331.38 ;
     RECT  210.61 252.88 217.79 331.38 ;
     RECT  300.21 264.88 307.39 331.38 ;
     RECT  379.54 329.7 396.99 331.38 ;
     RECT  793.01 252.88 800.19 331.38 ;
     RECT  823.06 330.63 823.34 331.38 ;
     RECT  837.81 252.88 844.99 331.38 ;
     RECT  379.54 331.38 410.62 331.66 ;
     RECT  524.21 252.88 550.62 331.66 ;
     RECT  160.02 328.39 176.54 333.62 ;
     RECT  191.38 331.38 191.66 333.62 ;
     RECT  255.41 252.88 262.59 333.62 ;
     RECT  327.46 330.82 352.19 333.62 ;
     RECT  454.02 330.82 463.26 333.62 ;
     RECT  927.41 252.88 934.59 333.62 ;
     RECT  296.66 331.38 307.39 334.18 ;
     RECT  919.94 333.62 934.59 334.18 ;
     RECT  703.41 252.88 710.59 334.74 ;
     RECT  722.26 334.18 722.54 334.74 ;
     RECT  917.7 334.18 934.59 334.74 ;
     RECT  524.21 331.66 549.5 335.58 ;
     RECT  76.21 252.88 83.39 336.42 ;
     RECT  379.54 331.66 396.99 336.42 ;
     RECT  453.46 333.62 463.26 336.42 ;
     RECT  602.98 330.26 620.99 336.42 ;
     RECT  453.46 336.42 464.38 338.38 ;
     RECT  9.94 328.39 38.59 339.78 ;
     RECT  658.61 252.88 665.79 340.9 ;
     RECT  972.21 330.82 991.34 340.9 ;
     RECT  434.61 252.88 441.79 341.46 ;
     RECT  972.21 340.9 993.02 342.146 ;
     RECT  858.9 341.46 859.18 343.98 ;
     RECT  972.21 342.146 1001.23 343.98 ;
     RECT  966.085 343.98 1001.23 344.26 ;
     RECT  965.3 344.26 1001.23 345.38 ;
     RECT  9.94 339.78 39.34 346.09 ;
     RECT  569.01 252.88 576.19 346.09 ;
     RECT  965.3 345.38 1004.22 348.18 ;
     RECT  565.74 346.09 576.19 348.74 ;
     RECT  858.9 343.98 863.885 349.3 ;
     RECT  965.3 348.18 1005.9 349.3 ;
     RECT  910.42 334.74 934.59 349.67 ;
     RECT  564.34 348.74 576.19 350.42 ;
     RECT  965.3 349.3 1006.46 350.495 ;
     RECT  429.94 341.46 441.79 350.98 ;
     RECT  454.02 338.38 464.38 350.98 ;
     RECT  910.42 349.67 940.94 350.98 ;
     RECT  9.94 346.09 42.42 352 ;
     RECT  76.21 336.42 91.42 352 ;
     RECT  121.01 331.38 140.14 352 ;
     RECT  160.02 333.62 191.66 352 ;
     RECT  210.61 331.38 223.58 352 ;
     RECT  255.41 333.62 272.3 352 ;
     RECT  292.74 334.18 307.39 352 ;
     RECT  326.9 333.62 352.19 352 ;
     RECT  376.18 336.42 396.99 352 ;
     RECT  429.94 350.98 464.38 352 ;
     RECT  524.21 335.58 545.58 352 ;
     RECT  560.42 350.42 576.19 352 ;
     RECT  602.98 336.42 622.3 352 ;
     RECT  658.61 340.9 671.02 352 ;
     RECT  690.9 333.62 691.18 352 ;
     RECT  703.41 334.74 722.54 352 ;
     RECT  748.21 330.63 764.54 352 ;
     RECT  793.01 331.38 803.18 352 ;
     RECT  823.06 331.38 844.99 352 ;
     RECT  858.9 349.3 866.74 352 ;
     RECT  882.61 252.88 889.79 352 ;
     RECT  907.06 350.98 940.94 352 ;
     RECT  961.1 350.495 1006.46 352 ;
     RECT  524.21 352 1006.46 355.74 ;
     RECT  9.94 352 464.38 357.98 ;
     RECT  524.21 355.74 1005.9 374.22 ;
     RECT  11.25 357.98 464.38 584.88 ;
     RECT  524.21 374.22 1001.23 584.88 ;
     RECT  11.25 584.88 16.19 590.254 ;
     RECT  993.49 584.88 1001.23 590.254 ;
     RECT  14.05 590.254 16.19 595.294 ;
     RECT  999.09 590.254 1001.23 595.294 ;
     RECT  434.61 584.88 464.38 596.26 ;
     RECT  604.66 584.88 626.78 596.54 ;
     RECT  429.94 596.26 464.38 598.22 ;
     RECT  524.21 584.88 545.58 598.22 ;
     RECT  385.7 584.88 396.99 598.5 ;
     RECT  429.94 598.22 454.3 598.78 ;
     RECT  545.3 598.22 545.58 598.78 ;
     RECT  376.18 598.5 396.99 599.62 ;
     RECT  610.82 596.54 626.78 601.58 ;
     RECT  375.9 599.62 396.99 602.57 ;
     RECT  429.94 598.78 452.62 603.54 ;
     RECT  31.41 584.88 38.59 605.374 ;
     RECT  76.21 584.88 83.39 605.374 ;
     RECT  121.01 584.88 128.19 605.374 ;
     RECT  165.81 584.88 172.99 605.374 ;
     RECT  210.61 584.88 217.79 605.374 ;
     RECT  255.41 584.88 262.59 605.374 ;
     RECT  300.21 584.88 307.39 605.374 ;
     RECT  345.01 584.88 352.19 605.374 ;
     RECT  479.41 192.78 486.59 605.374 ;
     RECT  524.21 598.22 531.39 605.374 ;
     RECT  658.61 584.88 665.79 605.374 ;
     RECT  703.41 584.88 710.59 605.374 ;
     RECT  748.21 584.88 755.39 605.374 ;
     RECT  793.01 584.88 800.19 605.374 ;
     RECT  837.81 584.88 844.99 605.374 ;
     RECT  882.61 584.88 889.79 605.374 ;
     RECT  927.41 584.88 934.59 605.374 ;
     RECT  972.21 584.88 979.39 605.374 ;
     RECT  410.9 584.88 411.18 606.06 ;
     RECT  429.66 603.54 452.62 606.9 ;
     RECT  610.82 601.58 629.02 606.9 ;
     RECT  567.14 584.88 576.19 607.03 ;
     RECT  435.54 606.9 452.62 607.18 ;
     RECT  561.26 607.03 576.19 607.74 ;
     RECT  379.54 602.57 396.99 608.02 ;
     RECT  435.54 607.18 445.34 608.02 ;
     RECT  561.26 607.74 576.94 608.02 ;
     RECT  616.98 606.9 629.02 608.86 ;
     RECT  561.26 608.02 561.54 610.26 ;
     RECT  36.45 605.374 38.59 610.414 ;
     RECT  81.25 605.374 83.39 610.414 ;
     RECT  126.05 605.374 128.19 610.414 ;
     RECT  170.85 605.374 172.99 610.414 ;
     RECT  215.65 605.374 217.79 610.414 ;
     RECT  260.45 605.374 262.59 610.414 ;
     RECT  305.25 605.374 307.39 610.414 ;
     RECT  350.05 605.374 352.19 610.414 ;
     RECT  392.98 608.02 396.99 610.414 ;
     RECT  435.54 608.02 441.79 610.414 ;
     RECT  484.45 605.374 486.59 610.414 ;
     RECT  529.25 605.374 531.39 610.414 ;
     RECT  574.05 608.02 576.94 610.414 ;
     RECT  618.85 608.86 629.02 610.414 ;
     RECT  663.65 605.374 665.79 610.414 ;
     RECT  708.45 605.374 710.59 610.414 ;
     RECT  753.25 605.374 755.39 610.414 ;
     RECT  798.05 605.374 800.19 610.414 ;
     RECT  842.85 605.374 844.99 610.414 ;
     RECT  887.65 605.374 889.79 610.414 ;
     RECT  932.45 605.374 934.59 610.414 ;
     RECT  977.25 605.374 979.39 610.414 ;
     RECT  379.54 608.02 380.1 610.54 ;
     RECT  560.98 610.26 561.54 610.54 ;
     RECT  620.9 610.414 629.02 611.66 ;
     RECT  379.54 610.54 379.82 612.78 ;
     RECT  435.54 610.414 439.18 612.78 ;
     RECT  560.98 610.54 561.26 612.78 ;
     RECT  392.98 610.414 393.82 613.34 ;
     RECT  435.54 612.78 435.82 613.34 ;
     RECT  576.1 610.414 576.94 613.34 ;
     RECT  620.9 611.66 621.74 613.9 ;
    LAYER Metal3 ;
     RECT  0.12 344.82 0.26 347.34 ;
     RECT  0.26 19.46 9.94 20.86 ;
     RECT  0.26 344.82 9.94 357.98 ;
     RECT  9.94 333.62 11.62 357.98 ;
     RECT  9.94 16.1 11.874 20.86 ;
     RECT  11.62 328.58 11.874 357.98 ;
     RECT  11.874 14.596 14.674 257.564 ;
     RECT  11.874 328.58 14.674 590.204 ;
     RECT  14.674 9.556 15.746 262.604 ;
     RECT  14.674 328.58 15.746 595.244 ;
     RECT  15.746 328.58 18.76 584.88 ;
     RECT  18.76 325.78 19.18 584.88 ;
     RECT  15.746 16.1 31.954 252.88 ;
     RECT  19.18 328.58 31.954 584.88 ;
     RECT  31.954 9.556 32.926 605.324 ;
     RECT  32.926 14.596 37.074 605.324 ;
     RECT  37.074 14.596 38.246 610.364 ;
     RECT  38.246 16.1 68.74 252.88 ;
     RECT  68.74 7.14 75.74 252.88 ;
     RECT  75.74 8.26 76.834 252.88 ;
     RECT  38.246 331.38 76.834 333.9 ;
     RECT  38.246 352 76.834 584.88 ;
     RECT  76.834 8.26 79.34 605.324 ;
     RECT  79.34 9.38 81.454 605.324 ;
     RECT  81.454 9.38 82.766 610.364 ;
     RECT  82.766 9.38 87.44 252.88 ;
     RECT  87.44 16.1 121.634 252.88 ;
     RECT  82.766 331.38 121.634 333.9 ;
     RECT  82.766 352 121.634 584.88 ;
     RECT  121.634 9.556 122.846 605.324 ;
     RECT  122.846 12.18 126.454 605.324 ;
     RECT  126.454 12.18 127.566 610.364 ;
     RECT  127.566 12.18 139.36 252.88 ;
     RECT  139.36 9.38 140.42 252.88 ;
     RECT  140.42 16.1 166.054 252.88 ;
     RECT  127.566 331.38 166.054 333.9 ;
     RECT  127.566 352 166.054 584.88 ;
     RECT  166.054 9.556 171.454 605.324 ;
     RECT  171.454 9.556 172.366 610.364 ;
     RECT  172.366 9.556 176.07 252.88 ;
     RECT  176.07 8.26 176.4 252.88 ;
     RECT  172.366 328.58 183.26 333.9 ;
     RECT  183.26 328.58 191.66 331.66 ;
     RECT  176.4 8.82 211.054 252.88 ;
     RECT  191.66 328.58 211.054 330.54 ;
     RECT  172.366 352 211.054 584.88 ;
     RECT  211.054 8.82 216.274 605.324 ;
     RECT  216.274 8.82 217.346 610.364 ;
     RECT  217.346 8.82 223.3 252.88 ;
     RECT  217.346 328.58 235.34 331.66 ;
     RECT  223.3 6.58 256.034 252.88 ;
     RECT  235.34 331.38 256.034 331.66 ;
     RECT  217.346 352 256.034 584.88 ;
     RECT  256.034 6.58 261.074 605.324 ;
     RECT  261.074 6.58 262.346 610.364 ;
     RECT  262.346 331.38 292.74 333.9 ;
     RECT  262.346 6.58 300.834 252.88 ;
     RECT  293.86 264.74 300.834 265.02 ;
     RECT  292.74 331.38 300.834 334.46 ;
     RECT  262.346 352 300.834 584.88 ;
     RECT  300.834 6.58 305.554 605.324 ;
     RECT  305.554 6.58 306.766 610.364 ;
     RECT  306.766 6.58 345.634 252.88 ;
     RECT  306.766 264.74 345.634 265.02 ;
     RECT  306.766 331.38 345.634 334.46 ;
     RECT  306.766 352 345.634 584.88 ;
     RECT  345.634 6.58 350.554 605.324 ;
     RECT  350.554 6.58 351.566 610.364 ;
     RECT  351.566 264.74 352.94 265.02 ;
     RECT  375.16 601.86 378.76 602.14 ;
     RECT  351.566 331.38 379.54 334.46 ;
     RECT  378.76 601.86 389.56 612.78 ;
     RECT  351.566 6.58 390.154 252.88 ;
     RECT  379.54 329.7 390.154 334.46 ;
     RECT  351.566 352 390.154 584.88 ;
     RECT  389.56 601.86 390.154 613.34 ;
     RECT  390.154 6.58 393.26 613.34 ;
     RECT  393.26 6.58 394.94 610.364 ;
     RECT  394.94 7.7 396.446 610.364 ;
     RECT  396.446 605.78 411.18 606.06 ;
     RECT  396.446 329.7 411.74 334.46 ;
     RECT  396.446 7.7 429.16 252.88 ;
     RECT  429.16 6.58 433.58 252.88 ;
     RECT  433.58 7.7 435.154 252.88 ;
     RECT  411.74 331.38 435.154 334.46 ;
     RECT  396.446 352 435.154 584.88 ;
     RECT  429.16 613.06 435.154 613.34 ;
     RECT  435.154 7.7 435.82 613.34 ;
     RECT  435.82 7.7 439.18 612.78 ;
     RECT  439.18 7.7 441.446 610.364 ;
     RECT  441.446 7.7 451.86 252.88 ;
     RECT  441.446 350.98 451.86 584.88 ;
     RECT  451.86 350.98 452.06 351.26 ;
     RECT  451.86 41.3 453.74 42.7 ;
     RECT  453.46 276.5 454.02 276.78 ;
     RECT  451.86 217.14 455.42 219.1 ;
     RECT  454.02 276.5 455.42 277.34 ;
     RECT  453.74 41.3 455.98 41.58 ;
     RECT  455.42 277.06 455.98 277.34 ;
     RECT  441.446 331.38 455.98 334.46 ;
     RECT  451.86 7.7 457.66 19.18 ;
     RECT  455.98 331.38 462.14 333.9 ;
     RECT  462.14 331.38 462.7 331.66 ;
     RECT  457.66 7.7 463.82 16.38 ;
     RECT  463.82 8.82 480.034 16.38 ;
     RECT  480.034 8.82 484.654 605.324 ;
     RECT  484.654 8.82 485.966 610.364 ;
     RECT  485.966 8.82 524.834 16.38 ;
     RECT  524.834 8.82 529.654 605.324 ;
     RECT  529.654 8.82 530.766 610.364 ;
     RECT  530.766 8.82 536.34 16.38 ;
     RECT  530.766 334.18 543.06 334.46 ;
     RECT  530.766 350.42 544.18 350.7 ;
     RECT  543.06 333.62 548.1 334.46 ;
     RECT  548.1 333.62 549.22 335.02 ;
     RECT  549.22 333.62 550.34 335.58 ;
     RECT  536.34 7.7 551 16.38 ;
     RECT  544.18 350.42 551 351.26 ;
     RECT  560.56 612.5 567.76 612.78 ;
     RECT  551 7.7 569.254 252.88 ;
     RECT  550.34 331.38 569.254 335.58 ;
     RECT  551 350.42 569.254 584.88 ;
     RECT  567.76 612.5 569.254 613.34 ;
     RECT  569.254 7.7 575.566 613.34 ;
     RECT  575.566 613.06 576.38 613.34 ;
     RECT  609.16 608.58 612.76 608.86 ;
     RECT  575.566 7.7 614.254 252.88 ;
     RECT  575.566 331.38 614.254 335.58 ;
     RECT  575.566 352 614.254 584.88 ;
     RECT  612.76 606.34 614.254 608.86 ;
     RECT  614.254 7.7 618.16 608.86 ;
     RECT  618.16 7.7 620.546 613.9 ;
     RECT  620.546 611.38 621.18 613.9 ;
     RECT  621.18 611.38 629.02 611.66 ;
     RECT  620.546 7.7 659.234 252.88 ;
     RECT  620.546 331.38 659.234 335.58 ;
     RECT  620.546 352 659.234 584.88 ;
     RECT  659.234 7.7 664.274 605.324 ;
     RECT  664.274 7.7 665.546 610.364 ;
     RECT  665.546 7.7 704.034 252.88 ;
     RECT  665.546 331.38 704.034 335.58 ;
     RECT  665.546 352 704.034 584.88 ;
     RECT  704.034 7.7 708.754 605.324 ;
     RECT  708.754 7.7 709.966 610.364 ;
     RECT  709.966 331.38 714.14 335.02 ;
     RECT  714.14 331.38 722.54 334.46 ;
     RECT  709.966 7.7 748.834 252.88 ;
     RECT  722.54 331.38 748.834 333.9 ;
     RECT  709.966 352 748.834 584.88 ;
     RECT  748.834 7.7 752.78 605.324 ;
     RECT  752.78 13.3 753.754 605.324 ;
     RECT  753.754 13.3 754.766 610.364 ;
     RECT  754.766 13.3 793.354 252.88 ;
     RECT  754.766 330.82 793.354 584.88 ;
     RECT  793.354 9.556 794.526 605.324 ;
     RECT  794.526 13.3 798.674 605.324 ;
     RECT  798.674 13.3 799.646 610.364 ;
     RECT  799.646 330.82 823.34 584.88 ;
     RECT  799.646 13.3 838.354 252.88 ;
     RECT  823.34 331.38 838.354 333.9 ;
     RECT  823.34 352 838.354 584.88 ;
     RECT  838.354 9.556 839.326 605.324 ;
     RECT  839.326 13.3 843.474 605.324 ;
     RECT  843.474 13.3 844.646 610.364 ;
     RECT  844.646 13.3 859.36 252.88 ;
     RECT  859.36 9.38 860.58 252.88 ;
     RECT  860.58 13.3 883.234 252.88 ;
     RECT  844.646 331.38 883.234 333.9 ;
     RECT  844.646 352 883.234 584.88 ;
     RECT  883.234 9.556 884.246 605.324 ;
     RECT  884.246 13.3 887.854 605.324 ;
     RECT  887.854 13.3 889.166 610.364 ;
     RECT  889.166 13.3 906.16 252.88 ;
     RECT  906.16 8.82 906.78 252.88 ;
     RECT  906.78 11.62 920.56 252.88 ;
     RECT  920.56 8.82 924.14 252.88 ;
     RECT  924.14 9.556 928.034 252.88 ;
     RECT  889.166 331.38 928.034 333.9 ;
     RECT  889.166 352 928.034 584.88 ;
     RECT  928.034 9.556 929.246 605.324 ;
     RECT  929.246 11.62 932.854 605.324 ;
     RECT  932.854 11.62 933.966 610.364 ;
     RECT  933.966 11.62 938.98 252.88 ;
     RECT  938.98 13.3 960.16 252.88 ;
     RECT  960.16 8.26 960.63 252.88 ;
     RECT  960.63 9.38 970.9 252.88 ;
     RECT  970.9 9.556 972.454 252.88 ;
     RECT  933.966 331.38 972.454 333.9 ;
     RECT  933.966 349.86 972.454 584.88 ;
     RECT  972.454 9.556 973.726 605.324 ;
     RECT  973.726 13.3 977.854 605.324 ;
     RECT  977.854 13.3 978.766 610.364 ;
     RECT  978.766 13.3 983.5 252.88 ;
     RECT  978.766 331.38 983.5 333.9 ;
     RECT  983.5 13.86 984.06 252.88 ;
     RECT  983.5 333.62 984.06 333.9 ;
     RECT  984.06 14.596 994.054 252.88 ;
     RECT  978.766 349.86 994.054 584.88 ;
     RECT  994.054 347.236 996.66 590.204 ;
     RECT  994.054 14.596 999.454 257.564 ;
     RECT  996.66 345.38 999.454 590.204 ;
     RECT  999.454 9.556 1000.606 262.604 ;
     RECT  999.454 342.196 1000.606 595.244 ;
     RECT  1000.606 345.38 1004.22 366.38 ;
     RECT  1004.22 347.62 1005.9 366.38 ;
     RECT  1005.9 347.62 1019.7 357.98 ;
    LAYER Metal4 ;
     RECT  75.38 0.9 81.22 1.12 ;
     RECT  390.38 0.9 394.42 1.12 ;
     RECT  568.58 0.9 570.82 1.12 ;
     RECT  618.98 0.9 623.92 1.12 ;
     RECT  910.58 0.9 920.02 1.12 ;
     RECT  429.08 1.12 438.52 5.94 ;
     RECT  429.08 5.94 439.42 6.94 ;
     RECT  609.08 1.12 623.92 8.06 ;
     RECT  160.88 1.12 175.72 8.18 ;
     RECT  160.88 8.18 176.62 8.62 ;
     RECT  609.08 8.06 622.16 8.62 ;
     RECT  960.08 1.12 969.52 8.62 ;
     RECT  906.08 1.12 920.92 9.18 ;
     RECT  75.38 1.12 91.12 9.506 ;
     RECT  132.08 1.12 139.72 9.506 ;
     RECT  328.28 1.12 335.92 9.506 ;
     RECT  360.68 1.12 394.42 9.506 ;
     RECT  488.48 1.12 488.92 9.506 ;
     RECT  560.48 1.12 570.82 9.506 ;
     RECT  663.08 1.12 670.72 9.506 ;
     RECT  859.28 1.12 866.92 9.506 ;
     RECT  915.08 9.18 920.92 9.506 ;
     RECT  969.08 8.62 969.52 9.506 ;
     RECT  119.84 9.506 139.72 9.74 ;
     RECT  328.28 9.506 394.42 9.74 ;
     RECT  560.48 9.506 572.32 9.74 ;
     RECT  859.28 9.506 885.92 9.74 ;
     RECT  969.08 9.506 975.52 9.74 ;
     RECT  657.44 9.506 670.72 11.54 ;
     RECT  657.44 11.54 671.62 11.98 ;
     RECT  915.08 9.506 930.72 11.98 ;
     RECT  119.84 9.74 132.52 12.54 ;
     RECT  478.24 9.506 488.92 12.54 ;
     RECT  919.58 11.98 930.72 12.54 ;
     RECT  335.48 9.74 370.12 13.66 ;
     RECT  14.18 9.506 34.72 14.546 ;
     RECT  209.44 9.506 213.92 14.546 ;
     RECT  254.24 9.506 258.72 14.546 ;
     RECT  299.04 9.506 303.52 14.546 ;
     RECT  388.64 9.74 394.42 14.546 ;
     RECT  433.44 6.94 439.42 14.546 ;
     RECT  523.04 9.506 527.52 14.546 ;
     RECT  567.84 9.74 572.32 14.546 ;
     RECT  702.24 9.506 706.72 14.546 ;
     RECT  747.04 9.506 751.52 14.546 ;
     RECT  791.84 9.506 796.32 14.546 ;
     RECT  836.64 9.506 841.12 14.546 ;
     RECT  866.48 9.74 885.92 14.546 ;
     RECT  926.24 12.54 930.72 14.546 ;
     RECT  971.04 9.74 975.52 14.546 ;
     RECT  997.66 9.506 1002.14 14.546 ;
     RECT  75.04 9.506 91.12 17.02 ;
     RECT  343.84 13.66 370.12 17.02 ;
     RECT  866.48 14.546 890.96 17.02 ;
     RECT  343.84 17.02 368.32 17.58 ;
     RECT  343.84 17.58 366.52 18.14 ;
     RECT  160.88 8.62 174.16 19.26 ;
     RECT  11.48 14.546 39.76 257.614 ;
     RECT  14.18 257.614 39.76 262.654 ;
     RECT  971.04 14.546 1002.14 262.654 ;
     RECT  30.24 262.654 39.76 325.7 ;
     RECT  18.68 325.7 39.76 342.146 ;
     RECT  971.04 262.654 980.56 342.146 ;
     RECT  14.18 342.146 39.76 347.186 ;
     RECT  11.48 347.186 39.76 590.254 ;
     RECT  14.18 590.254 39.76 595.294 ;
     RECT  971.04 342.146 1002.14 595.294 ;
     RECT  388.64 14.546 398.16 601.78 ;
     RECT  30.24 595.294 39.76 605.374 ;
     RECT  75.04 17.02 84.56 605.374 ;
     RECT  119.84 12.54 129.36 605.374 ;
     RECT  164.64 19.26 174.16 605.374 ;
     RECT  209.44 14.546 218.96 605.374 ;
     RECT  254.24 14.546 263.76 605.374 ;
     RECT  299.04 14.546 308.56 605.374 ;
     RECT  343.84 18.14 353.36 605.374 ;
     RECT  478.24 12.54 487.76 605.374 ;
     RECT  523.04 14.546 532.56 605.374 ;
     RECT  657.44 11.98 666.96 605.374 ;
     RECT  702.24 14.546 711.76 605.374 ;
     RECT  747.04 14.546 756.56 605.374 ;
     RECT  791.84 14.546 801.36 605.374 ;
     RECT  836.64 14.546 846.16 605.374 ;
     RECT  881.44 17.02 890.96 605.374 ;
     RECT  926.24 14.546 935.76 605.374 ;
     RECT  971.04 595.294 980.56 605.374 ;
     RECT  612.64 8.62 622.16 608.5 ;
     RECT  35.28 605.374 39.76 610.414 ;
     RECT  80.08 605.374 84.56 610.414 ;
     RECT  124.88 605.374 129.36 610.414 ;
     RECT  169.68 605.374 174.16 610.414 ;
     RECT  214.48 605.374 218.96 610.414 ;
     RECT  259.28 605.374 263.76 610.414 ;
     RECT  304.08 605.374 308.56 610.414 ;
     RECT  348.88 605.374 353.36 610.414 ;
     RECT  375.08 601.78 398.16 610.414 ;
     RECT  433.44 14.546 442.96 610.414 ;
     RECT  483.28 605.374 487.76 610.414 ;
     RECT  528.08 605.374 532.56 610.414 ;
     RECT  567.84 14.546 577.36 610.414 ;
     RECT  609.08 608.5 622.16 610.414 ;
     RECT  662.48 605.374 666.96 610.414 ;
     RECT  707.28 605.374 711.76 610.414 ;
     RECT  752.08 605.374 756.56 610.414 ;
     RECT  796.88 605.374 801.36 610.414 ;
     RECT  841.68 605.374 846.16 610.414 ;
     RECT  886.48 605.374 890.96 610.414 ;
     RECT  931.28 605.374 935.76 610.414 ;
     RECT  976.08 605.374 980.56 610.414 ;
     RECT  567.84 610.414 568.12 612.42 ;
     RECT  433.44 610.414 438.52 612.98 ;
     RECT  375.08 610.414 389.92 618.8 ;
     RECT  429.08 612.98 438.52 618.8 ;
     RECT  560.48 612.42 568.12 618.8 ;
     RECT  609.08 610.414 622.12 618.8 ;
  END
END mem_64_32_gf180
END LIBRARY
