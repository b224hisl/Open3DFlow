VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO mem_64_16_gf180
  FOREIGN mem_64_16_gf180 0 0 ;
  CLASS BLOCK ;
  SIZE 620 BY 610.414 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  572.88 14.546 577.36 610.414 ;
        RECT  528.08 14.546 532.56 610.414 ;
        RECT  483.28 14.546 487.76 610.414 ;
        RECT  438.48 14.546 442.96 610.414 ;
        RECT  393.68 14.546 398.16 610.414 ;
        RECT  348.88 14.546 353.36 610.414 ;
        RECT  304.08 14.546 308.56 610.414 ;
        RECT  259.28 14.546 263.76 610.414 ;
        RECT  214.48 14.546 218.96 610.414 ;
        RECT  169.68 14.546 174.16 610.414 ;
        RECT  124.88 14.546 129.36 610.414 ;
        RECT  80.08 14.546 84.56 610.414 ;
        RECT  35.28 14.546 39.76 610.414 ;
      LAYER Metal1 ;
        RECT  528.08 599.31 609.84 600.21 ;
        RECT  528.08 589.23 609.84 590.13 ;
        RECT  528.08 579.15 609.84 580.05 ;
        RECT  528.08 569.07 609.84 569.97 ;
        RECT  528.08 558.99 609.84 559.89 ;
        RECT  528.08 548.91 609.84 549.81 ;
        RECT  528.08 538.83 609.84 539.73 ;
        RECT  528.08 528.75 609.84 529.65 ;
        RECT  528.08 518.67 609.84 519.57 ;
        RECT  528.08 508.59 609.84 509.49 ;
        RECT  528.08 498.51 609.84 499.41 ;
        RECT  528.08 488.43 609.84 489.33 ;
        RECT  528.08 478.35 609.84 479.25 ;
        RECT  528.08 468.27 609.84 469.17 ;
        RECT  528.08 458.19 609.84 459.09 ;
        RECT  528.08 448.11 609.84 449.01 ;
        RECT  528.08 438.03 609.84 438.93 ;
        RECT  528.08 427.95 609.84 428.85 ;
        RECT  528.08 417.87 609.84 418.77 ;
        RECT  528.08 407.79 609.84 408.69 ;
        RECT  528.08 397.71 609.84 398.61 ;
        RECT  528.08 387.63 609.84 388.53 ;
        RECT  528.08 377.55 609.84 378.45 ;
        RECT  528.08 367.47 609.84 368.37 ;
        RECT  528.08 246.51 609.84 247.41 ;
        RECT  528.08 236.43 609.84 237.33 ;
        RECT  528.08 226.35 609.84 227.25 ;
        RECT  528.08 216.27 609.84 217.17 ;
        RECT  528.08 206.19 609.84 207.09 ;
        RECT  528.08 196.11 609.84 197.01 ;
        RECT  528.08 186.03 609.84 186.93 ;
        RECT  528.08 175.95 609.84 176.85 ;
        RECT  528.08 165.87 609.84 166.77 ;
        RECT  528.08 155.79 609.84 156.69 ;
        RECT  528.08 145.71 609.84 146.61 ;
        RECT  528.08 135.63 609.84 136.53 ;
        RECT  528.08 125.55 609.84 126.45 ;
        RECT  528.08 115.47 609.84 116.37 ;
        RECT  528.08 105.39 609.84 106.29 ;
        RECT  528.08 95.31 609.84 96.21 ;
        RECT  528.08 85.23 609.84 86.13 ;
        RECT  528.08 75.15 609.84 76.05 ;
        RECT  528.08 65.07 609.84 65.97 ;
        RECT  528.08 54.99 609.84 55.89 ;
        RECT  528.08 44.91 609.84 45.81 ;
        RECT  528.08 34.83 609.84 35.73 ;
        RECT  528.08 24.75 609.84 25.65 ;
        RECT  10.08 609.39 609.84 610.29 ;
        RECT  10.08 599.31 92.96 600.21 ;
        RECT  10.08 589.23 92.96 590.13 ;
        RECT  10.08 579.15 92.96 580.05 ;
        RECT  10.08 569.07 92.96 569.97 ;
        RECT  10.08 558.99 92.96 559.89 ;
        RECT  10.08 548.91 92.96 549.81 ;
        RECT  10.08 538.83 92.96 539.73 ;
        RECT  10.08 528.75 92.96 529.65 ;
        RECT  10.08 518.67 92.96 519.57 ;
        RECT  10.08 508.59 92.96 509.49 ;
        RECT  10.08 498.51 92.96 499.41 ;
        RECT  10.08 488.43 92.96 489.33 ;
        RECT  10.08 478.35 92.96 479.25 ;
        RECT  10.08 468.27 92.96 469.17 ;
        RECT  10.08 458.19 92.96 459.09 ;
        RECT  10.08 448.11 92.96 449.01 ;
        RECT  10.08 438.03 92.96 438.93 ;
        RECT  10.08 427.95 92.96 428.85 ;
        RECT  10.08 417.87 92.96 418.77 ;
        RECT  10.08 407.79 92.96 408.69 ;
        RECT  10.08 397.71 92.96 398.61 ;
        RECT  10.08 387.63 92.96 388.53 ;
        RECT  10.08 377.55 92.96 378.45 ;
        RECT  10.08 367.47 92.96 368.37 ;
        RECT  10.08 357.39 609.84 358.29 ;
        RECT  10.08 347.31 609.84 348.21 ;
        RECT  10.08 337.23 609.84 338.13 ;
        RECT  10.08 327.15 609.84 328.05 ;
        RECT  10.08 317.07 609.84 317.97 ;
        RECT  10.08 306.99 609.84 307.89 ;
        RECT  10.08 296.91 609.84 297.81 ;
        RECT  10.08 286.83 609.84 287.73 ;
        RECT  10.08 276.75 609.84 277.65 ;
        RECT  10.08 266.67 609.84 267.57 ;
        RECT  10.08 256.59 609.84 257.49 ;
        RECT  10.08 246.51 92.96 247.41 ;
        RECT  10.08 236.43 92.96 237.33 ;
        RECT  10.08 226.35 92.96 227.25 ;
        RECT  10.08 216.27 92.96 217.17 ;
        RECT  10.08 206.19 92.96 207.09 ;
        RECT  10.08 196.11 92.96 197.01 ;
        RECT  10.08 186.03 92.96 186.93 ;
        RECT  10.08 175.95 92.96 176.85 ;
        RECT  10.08 165.87 92.96 166.77 ;
        RECT  10.08 155.79 92.96 156.69 ;
        RECT  10.08 145.71 92.96 146.61 ;
        RECT  10.08 135.63 92.96 136.53 ;
        RECT  10.08 125.55 92.96 126.45 ;
        RECT  10.08 115.47 92.96 116.37 ;
        RECT  10.08 105.39 92.96 106.29 ;
        RECT  10.08 95.31 92.96 96.21 ;
        RECT  10.08 85.23 92.96 86.13 ;
        RECT  10.08 75.15 92.96 76.05 ;
        RECT  10.08 65.07 92.96 65.97 ;
        RECT  10.08 54.99 92.96 55.89 ;
        RECT  10.08 44.91 92.96 45.81 ;
        RECT  10.08 34.83 92.96 35.73 ;
        RECT  10.08 24.75 92.96 25.65 ;
        RECT  10.08 14.67 609.84 15.57 ;
      VIA 575.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 609.266 576.19 610.414 ;
      VIA 575.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 599.186 576.19 600.334 ;
      VIA 575.376 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 589.106 576.19 590.254 ;
      VIA 575.376 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 579.026 576.19 580.174 ;
      VIA 575.376 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 568.946 576.19 570.094 ;
      VIA 575.376 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 558.866 576.19 560.014 ;
      VIA 575.376 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 548.786 576.19 549.934 ;
      VIA 575.376 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 538.706 576.19 539.854 ;
      VIA 575.376 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 528.626 576.19 529.774 ;
      VIA 575.376 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 518.546 576.19 519.694 ;
      VIA 575.376 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 508.466 576.19 509.614 ;
      VIA 575.376 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 498.386 576.19 499.534 ;
      VIA 575.376 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 488.306 576.19 489.454 ;
      VIA 575.376 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 478.226 576.19 479.374 ;
      VIA 575.376 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 468.146 576.19 469.294 ;
      VIA 575.376 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 458.066 576.19 459.214 ;
      VIA 575.376 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 447.986 576.19 449.134 ;
      VIA 575.376 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 437.906 576.19 439.054 ;
      VIA 575.376 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 427.826 576.19 428.974 ;
      VIA 575.376 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 417.746 576.19 418.894 ;
      VIA 575.376 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 407.666 576.19 408.814 ;
      VIA 575.376 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 397.586 576.19 398.734 ;
      VIA 575.376 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 387.506 576.19 388.654 ;
      VIA 575.376 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 377.426 576.19 378.574 ;
      VIA 575.376 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 367.346 576.19 368.494 ;
      VIA 575.376 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 357.266 576.19 358.414 ;
      VIA 575.376 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 347.186 576.19 348.334 ;
      VIA 575.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 337.106 576.19 338.254 ;
      VIA 575.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 327.026 576.19 328.174 ;
      VIA 575.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 316.946 576.19 318.094 ;
      VIA 575.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 306.866 576.19 308.014 ;
      VIA 575.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 296.786 576.19 297.934 ;
      VIA 575.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 286.706 576.19 287.854 ;
      VIA 575.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 276.626 576.19 277.774 ;
      VIA 575.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 266.546 576.19 267.694 ;
      VIA 575.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 256.466 576.19 257.614 ;
      VIA 575.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 246.386 576.19 247.534 ;
      VIA 575.376 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 236.306 576.19 237.454 ;
      VIA 575.376 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 226.226 576.19 227.374 ;
      VIA 575.376 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 216.146 576.19 217.294 ;
      VIA 575.376 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 206.066 576.19 207.214 ;
      VIA 575.376 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 195.986 576.19 197.134 ;
      VIA 575.376 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 185.906 576.19 187.054 ;
      VIA 575.376 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 175.826 576.19 176.974 ;
      VIA 575.376 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 165.746 576.19 166.894 ;
      VIA 575.376 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 155.666 576.19 156.814 ;
      VIA 575.376 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 145.586 576.19 146.734 ;
      VIA 575.376 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 135.506 576.19 136.654 ;
      VIA 575.376 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 125.426 576.19 126.574 ;
      VIA 575.376 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 115.346 576.19 116.494 ;
      VIA 575.376 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 105.266 576.19 106.414 ;
      VIA 575.376 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 95.186 576.19 96.334 ;
      VIA 575.376 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 85.106 576.19 86.254 ;
      VIA 575.376 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 75.026 576.19 76.174 ;
      VIA 575.376 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 64.946 576.19 66.094 ;
      VIA 575.376 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 54.866 576.19 56.014 ;
      VIA 575.376 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 44.786 576.19 45.934 ;
      VIA 575.376 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 34.706 576.19 35.854 ;
      VIA 575.376 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 24.626 576.19 25.774 ;
      VIA 575.376 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 575.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 575.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 574.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  574.05 14.546 576.19 15.694 ;
      VIA 575.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 574.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 575.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 609.266 531.39 610.414 ;
      VIA 530.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 599.186 531.39 600.334 ;
      VIA 530.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 589.106 531.39 590.254 ;
      VIA 530.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 579.026 531.39 580.174 ;
      VIA 530.576 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 568.946 531.39 570.094 ;
      VIA 530.576 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 558.866 531.39 560.014 ;
      VIA 530.576 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 548.786 531.39 549.934 ;
      VIA 530.576 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 538.706 531.39 539.854 ;
      VIA 530.576 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 528.626 531.39 529.774 ;
      VIA 530.576 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 518.546 531.39 519.694 ;
      VIA 530.576 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 508.466 531.39 509.614 ;
      VIA 530.576 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 498.386 531.39 499.534 ;
      VIA 530.576 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 488.306 531.39 489.454 ;
      VIA 530.576 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 478.226 531.39 479.374 ;
      VIA 530.576 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 468.146 531.39 469.294 ;
      VIA 530.576 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 458.066 531.39 459.214 ;
      VIA 530.576 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 447.986 531.39 449.134 ;
      VIA 530.576 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 437.906 531.39 439.054 ;
      VIA 530.576 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 427.826 531.39 428.974 ;
      VIA 530.576 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 417.746 531.39 418.894 ;
      VIA 530.576 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 407.666 531.39 408.814 ;
      VIA 530.576 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 397.586 531.39 398.734 ;
      VIA 530.576 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 387.506 531.39 388.654 ;
      VIA 530.576 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 377.426 531.39 378.574 ;
      VIA 530.576 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 367.346 531.39 368.494 ;
      VIA 530.576 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 357.266 531.39 358.414 ;
      VIA 530.576 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 347.186 531.39 348.334 ;
      VIA 530.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 337.106 531.39 338.254 ;
      VIA 530.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 327.026 531.39 328.174 ;
      VIA 530.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 316.946 531.39 318.094 ;
      VIA 530.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 306.866 531.39 308.014 ;
      VIA 530.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 296.786 531.39 297.934 ;
      VIA 530.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 286.706 531.39 287.854 ;
      VIA 530.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 276.626 531.39 277.774 ;
      VIA 530.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 266.546 531.39 267.694 ;
      VIA 530.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 256.466 531.39 257.614 ;
      VIA 530.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 246.386 531.39 247.534 ;
      VIA 530.576 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 236.306 531.39 237.454 ;
      VIA 530.576 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 226.226 531.39 227.374 ;
      VIA 530.576 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 216.146 531.39 217.294 ;
      VIA 530.576 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 206.066 531.39 207.214 ;
      VIA 530.576 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 195.986 531.39 197.134 ;
      VIA 530.576 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 185.906 531.39 187.054 ;
      VIA 530.576 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 175.826 531.39 176.974 ;
      VIA 530.576 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 165.746 531.39 166.894 ;
      VIA 530.576 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 155.666 531.39 156.814 ;
      VIA 530.576 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 145.586 531.39 146.734 ;
      VIA 530.576 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 135.506 531.39 136.654 ;
      VIA 530.576 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 125.426 531.39 126.574 ;
      VIA 530.576 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 115.346 531.39 116.494 ;
      VIA 530.576 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 105.266 531.39 106.414 ;
      VIA 530.576 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 95.186 531.39 96.334 ;
      VIA 530.576 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 85.106 531.39 86.254 ;
      VIA 530.576 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 75.026 531.39 76.174 ;
      VIA 530.576 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 64.946 531.39 66.094 ;
      VIA 530.576 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 54.866 531.39 56.014 ;
      VIA 530.576 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 44.786 531.39 45.934 ;
      VIA 530.576 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 34.706 531.39 35.854 ;
      VIA 530.576 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 24.626 531.39 25.774 ;
      VIA 530.576 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 530.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 530.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 529.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  529.25 14.546 531.39 15.694 ;
      VIA 530.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 530.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 609.266 486.59 610.414 ;
      VIA 485.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 357.266 486.59 358.414 ;
      VIA 485.776 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 347.186 486.59 348.334 ;
      VIA 485.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 337.106 486.59 338.254 ;
      VIA 485.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 327.026 486.59 328.174 ;
      VIA 485.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 316.946 486.59 318.094 ;
      VIA 485.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 306.866 486.59 308.014 ;
      VIA 485.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 296.786 486.59 297.934 ;
      VIA 485.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 286.706 486.59 287.854 ;
      VIA 485.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 276.626 486.59 277.774 ;
      VIA 485.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 266.546 486.59 267.694 ;
      VIA 485.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 256.466 486.59 257.614 ;
      VIA 485.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 485.356 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.356 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.228 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 485.1 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.972 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 484.844 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  484.45 14.546 486.59 15.694 ;
      VIA 485.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 485.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 609.266 441.79 610.414 ;
      VIA 440.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 357.266 441.79 358.414 ;
      VIA 440.976 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 347.186 441.79 348.334 ;
      VIA 440.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 337.106 441.79 338.254 ;
      VIA 440.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 327.026 441.79 328.174 ;
      VIA 440.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 316.946 441.79 318.094 ;
      VIA 440.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 306.866 441.79 308.014 ;
      VIA 440.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 296.786 441.79 297.934 ;
      VIA 440.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 286.706 441.79 287.854 ;
      VIA 440.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 276.626 441.79 277.774 ;
      VIA 440.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 266.546 441.79 267.694 ;
      VIA 440.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 256.466 441.79 257.614 ;
      VIA 440.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 441.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 441 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 440.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  439.65 14.546 441.79 15.694 ;
      VIA 440.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 440.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 609.266 396.99 610.414 ;
      VIA 396.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 357.266 396.99 358.414 ;
      VIA 396.176 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 347.186 396.99 348.334 ;
      VIA 396.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 337.106 396.99 338.254 ;
      VIA 396.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 327.026 396.99 328.174 ;
      VIA 396.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 316.946 396.99 318.094 ;
      VIA 396.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 306.866 396.99 308.014 ;
      VIA 396.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 296.786 396.99 297.934 ;
      VIA 396.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 286.706 396.99 287.854 ;
      VIA 396.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 276.626 396.99 277.774 ;
      VIA 396.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 266.546 396.99 267.694 ;
      VIA 396.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 256.466 396.99 257.614 ;
      VIA 396.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 396.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 396 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 395.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  394.85 14.546 396.99 15.694 ;
      VIA 396.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 396.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 395.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 609.266 352.19 610.414 ;
      VIA 351.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 357.266 352.19 358.414 ;
      VIA 351.376 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 347.186 352.19 348.334 ;
      VIA 351.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 337.106 352.19 338.254 ;
      VIA 351.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 327.026 352.19 328.174 ;
      VIA 351.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 316.946 352.19 318.094 ;
      VIA 351.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 306.866 352.19 308.014 ;
      VIA 351.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 296.786 352.19 297.934 ;
      VIA 351.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 286.706 352.19 287.854 ;
      VIA 351.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 276.626 352.19 277.774 ;
      VIA 351.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 266.546 352.19 267.694 ;
      VIA 351.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 256.466 352.19 257.614 ;
      VIA 351.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 351.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 351 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 350.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  350.05 14.546 352.19 15.694 ;
      VIA 351.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 350.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 351.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 609.266 307.39 610.414 ;
      VIA 306.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 357.266 307.39 358.414 ;
      VIA 306.576 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 347.186 307.39 348.334 ;
      VIA 306.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 337.106 307.39 338.254 ;
      VIA 306.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 327.026 307.39 328.174 ;
      VIA 306.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 316.946 307.39 318.094 ;
      VIA 306.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 306.866 307.39 308.014 ;
      VIA 306.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 296.786 307.39 297.934 ;
      VIA 306.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 286.706 307.39 287.854 ;
      VIA 306.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 276.626 307.39 277.774 ;
      VIA 306.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 266.546 307.39 267.694 ;
      VIA 306.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 256.466 307.39 257.614 ;
      VIA 306.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 306.256 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.256 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306.128 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 306 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.872 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 305.744 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  305.25 14.546 307.39 15.694 ;
      VIA 306.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 306.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 609.266 262.59 610.414 ;
      VIA 261.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 357.266 262.59 358.414 ;
      VIA 261.776 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 347.186 262.59 348.334 ;
      VIA 261.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 337.106 262.59 338.254 ;
      VIA 261.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 327.026 262.59 328.174 ;
      VIA 261.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 316.946 262.59 318.094 ;
      VIA 261.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 306.866 262.59 308.014 ;
      VIA 261.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 296.786 262.59 297.934 ;
      VIA 261.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 286.706 262.59 287.854 ;
      VIA 261.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 276.626 262.59 277.774 ;
      VIA 261.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 266.546 262.59 267.694 ;
      VIA 261.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 256.466 262.59 257.614 ;
      VIA 261.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 262.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 262.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 261.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  260.45 14.546 262.59 15.694 ;
      VIA 261.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 261.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 609.266 217.79 610.414 ;
      VIA 216.976 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 357.266 217.79 358.414 ;
      VIA 216.976 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 347.186 217.79 348.334 ;
      VIA 216.976 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 337.106 217.79 338.254 ;
      VIA 216.976 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 327.026 217.79 328.174 ;
      VIA 216.976 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 316.946 217.79 318.094 ;
      VIA 216.976 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 306.866 217.79 308.014 ;
      VIA 216.976 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 296.786 217.79 297.934 ;
      VIA 216.976 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 286.706 217.79 287.854 ;
      VIA 216.976 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 276.626 217.79 277.774 ;
      VIA 216.976 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 266.546 217.79 267.694 ;
      VIA 216.976 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 256.466 217.79 257.614 ;
      VIA 216.976 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 217.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 217.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 216.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  215.65 14.546 217.79 15.694 ;
      VIA 216.976 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.976 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.848 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.592 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.464 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 216.72 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 609.266 172.99 610.414 ;
      VIA 172.176 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 357.266 172.99 358.414 ;
      VIA 172.176 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 347.186 172.99 348.334 ;
      VIA 172.176 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 337.106 172.99 338.254 ;
      VIA 172.176 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 327.026 172.99 328.174 ;
      VIA 172.176 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 316.946 172.99 318.094 ;
      VIA 172.176 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 306.866 172.99 308.014 ;
      VIA 172.176 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 296.786 172.99 297.934 ;
      VIA 172.176 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 286.706 172.99 287.854 ;
      VIA 172.176 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 276.626 172.99 277.774 ;
      VIA 172.176 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 266.546 172.99 267.694 ;
      VIA 172.176 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 256.466 172.99 257.614 ;
      VIA 172.176 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 172.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 172.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 171.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  170.85 14.546 172.99 15.694 ;
      VIA 172.176 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.176 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 172.048 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.792 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.664 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 171.92 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 609.266 128.19 610.414 ;
      VIA 127.376 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 357.266 128.19 358.414 ;
      VIA 127.376 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 347.186 128.19 348.334 ;
      VIA 127.376 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 337.106 128.19 338.254 ;
      VIA 127.376 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 327.026 128.19 328.174 ;
      VIA 127.376 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 316.946 128.19 318.094 ;
      VIA 127.376 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 306.866 128.19 308.014 ;
      VIA 127.376 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 296.786 128.19 297.934 ;
      VIA 127.376 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 286.706 128.19 287.854 ;
      VIA 127.376 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 276.626 128.19 277.774 ;
      VIA 127.376 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 266.546 128.19 267.694 ;
      VIA 127.376 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 256.466 128.19 257.614 ;
      VIA 127.376 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 127.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 127.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 126.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  126.05 14.546 128.19 15.694 ;
      VIA 127.376 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.376 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.248 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.992 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 126.864 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 127.12 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 609.266 83.39 610.414 ;
      VIA 82.576 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 599.186 83.39 600.334 ;
      VIA 82.576 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 589.106 83.39 590.254 ;
      VIA 82.576 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 579.026 83.39 580.174 ;
      VIA 82.576 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 568.946 83.39 570.094 ;
      VIA 82.576 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 558.866 83.39 560.014 ;
      VIA 82.576 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 548.786 83.39 549.934 ;
      VIA 82.576 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 538.706 83.39 539.854 ;
      VIA 82.576 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 528.626 83.39 529.774 ;
      VIA 82.576 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 518.546 83.39 519.694 ;
      VIA 82.576 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 508.466 83.39 509.614 ;
      VIA 82.576 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 498.386 83.39 499.534 ;
      VIA 82.576 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 488.306 83.39 489.454 ;
      VIA 82.576 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 478.226 83.39 479.374 ;
      VIA 82.576 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 468.146 83.39 469.294 ;
      VIA 82.576 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 458.066 83.39 459.214 ;
      VIA 82.576 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 447.986 83.39 449.134 ;
      VIA 82.576 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 437.906 83.39 439.054 ;
      VIA 82.576 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 427.826 83.39 428.974 ;
      VIA 82.576 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 417.746 83.39 418.894 ;
      VIA 82.576 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 407.666 83.39 408.814 ;
      VIA 82.576 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 397.586 83.39 398.734 ;
      VIA 82.576 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 387.506 83.39 388.654 ;
      VIA 82.576 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 377.426 83.39 378.574 ;
      VIA 82.576 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 367.346 83.39 368.494 ;
      VIA 82.576 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 357.266 83.39 358.414 ;
      VIA 82.576 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 347.186 83.39 348.334 ;
      VIA 82.576 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 337.106 83.39 338.254 ;
      VIA 82.576 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 327.026 83.39 328.174 ;
      VIA 82.576 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 316.946 83.39 318.094 ;
      VIA 82.576 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 306.866 83.39 308.014 ;
      VIA 82.576 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 296.786 83.39 297.934 ;
      VIA 82.576 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 286.706 83.39 287.854 ;
      VIA 82.576 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 276.626 83.39 277.774 ;
      VIA 82.576 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 266.546 83.39 267.694 ;
      VIA 82.576 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 256.466 83.39 257.614 ;
      VIA 82.576 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 246.386 83.39 247.534 ;
      VIA 82.576 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 236.306 83.39 237.454 ;
      VIA 82.576 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 226.226 83.39 227.374 ;
      VIA 82.576 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 216.146 83.39 217.294 ;
      VIA 82.576 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 206.066 83.39 207.214 ;
      VIA 82.576 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 195.986 83.39 197.134 ;
      VIA 82.576 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 185.906 83.39 187.054 ;
      VIA 82.576 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 175.826 83.39 176.974 ;
      VIA 82.576 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 165.746 83.39 166.894 ;
      VIA 82.576 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 155.666 83.39 156.814 ;
      VIA 82.576 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 145.586 83.39 146.734 ;
      VIA 82.576 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 135.506 83.39 136.654 ;
      VIA 82.576 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 125.426 83.39 126.574 ;
      VIA 82.576 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 115.346 83.39 116.494 ;
      VIA 82.576 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 105.266 83.39 106.414 ;
      VIA 82.576 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 95.186 83.39 96.334 ;
      VIA 82.576 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 85.106 83.39 86.254 ;
      VIA 82.576 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 75.026 83.39 76.174 ;
      VIA 82.576 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 64.946 83.39 66.094 ;
      VIA 82.576 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 54.866 83.39 56.014 ;
      VIA 82.576 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 44.786 83.39 45.934 ;
      VIA 82.576 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 34.706 83.39 35.854 ;
      VIA 82.576 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 24.626 83.39 25.774 ;
      VIA 82.576 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 82.156 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.156 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 82.028 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.9 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.772 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 81.644 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  81.25 14.546 83.39 15.694 ;
      VIA 82.576 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.576 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.448 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.192 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.064 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 82.32 15.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 610.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 610.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 609.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 609.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 609.266 38.59 610.414 ;
      VIA 37.776 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 610.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 610.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 609.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 609.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 600.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 600.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 599.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 599.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 599.186 38.59 600.334 ;
      VIA 37.776 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 600.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 600.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 599.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 599.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 590.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 589.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 589.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 589.106 38.59 590.254 ;
      VIA 37.776 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 590.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 589.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 589.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 579.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 579.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 579.026 38.59 580.174 ;
      VIA 37.776 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 579.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 579.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 569.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 569.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 568.946 38.59 570.094 ;
      VIA 37.776 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 569.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 569.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 559.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 559.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 558.866 38.59 560.014 ;
      VIA 37.776 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 559.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 559.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 549.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 548.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 548.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 548.786 38.59 549.934 ;
      VIA 37.776 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 549.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 548.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 549.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 539.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 538.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 538.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 538.706 38.59 539.854 ;
      VIA 37.776 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 539.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 538.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 539.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 529.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 529.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 529.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 529.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 529.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 528.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 528.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 528.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 528.626 38.59 529.774 ;
      VIA 37.776 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 529.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 529.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 529.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 529.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 529.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 528.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 528.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 529.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 519.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 519.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 519.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 519.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 518.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 518.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 518.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 518.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 518.546 38.59 519.694 ;
      VIA 37.776 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 519.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 519.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 519.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 519.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 518.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 518.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 518.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 519.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 509.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 509.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 509.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 509.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 508.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 508.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 508.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 508.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 508.466 38.59 509.614 ;
      VIA 37.776 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 509.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 509.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 509.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 509.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 508.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 508.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 508.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 509.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 499.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 499.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 499.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 498.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 498.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 498.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 498.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 498.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 498.386 38.59 499.534 ;
      VIA 37.776 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 499.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 499.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 499.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 498.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 498.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 498.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 498.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 498.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 489.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 489.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 489.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 488.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 488.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 488.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 488.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 488.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 488.306 38.59 489.454 ;
      VIA 37.776 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 489.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 489.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 489.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 488.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 488.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 488.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 488.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 488.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 479.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 479.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 478.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 478.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 478.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 478.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 478.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 478.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 478.226 38.59 479.374 ;
      VIA 37.776 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 479.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 479.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 478.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 478.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 478.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 478.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 478.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 478.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 469.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 468.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 468.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 468.146 38.59 469.294 ;
      VIA 37.776 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 469.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 468.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 468.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 459.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 458.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 458.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 458.066 38.59 459.214 ;
      VIA 37.776 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 459.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 458.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 458.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 448.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 448.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 447.986 38.59 449.134 ;
      VIA 37.776 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 448.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 448.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 438.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 438.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 437.906 38.59 439.054 ;
      VIA 37.776 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 438.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 438.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 428.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 428.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 427.826 38.59 428.974 ;
      VIA 37.776 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 428.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 428.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 418.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 417.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 417.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 417.746 38.59 418.894 ;
      VIA 37.776 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 418.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 417.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 418.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 408.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 408.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 408.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 408.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 408.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 407.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 407.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 407.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 407.666 38.59 408.814 ;
      VIA 37.776 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 408.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 408.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 408.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 408.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 408.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 407.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 407.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 408.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 398.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 398.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 398.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 398.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 398.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 397.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 397.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 397.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 397.586 38.59 398.734 ;
      VIA 37.776 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 398.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 398.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 398.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 398.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 398.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 397.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 397.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 398.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 388.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 388.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 388.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 388.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 387.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 387.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 387.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 387.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 387.506 38.59 388.654 ;
      VIA 37.776 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 388.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 388.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 388.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 388.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 387.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 387.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 387.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 388.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 378.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 378.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 378.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 378 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 377.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 377.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 377.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 377.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 377.426 38.59 378.574 ;
      VIA 37.776 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 378.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 378.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 378.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 378 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 377.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 377.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 377.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 378 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 368.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 368.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 368.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 367.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 367.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 367.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 367.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 367.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 367.346 38.59 368.494 ;
      VIA 37.776 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 368.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 368.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 368.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 367.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 367.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 367.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 367.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 367.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 358.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 358.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 357.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 357.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 357.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 357.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 357.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 357.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 357.266 38.59 358.414 ;
      VIA 37.776 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 358.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 358.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 357.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 357.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 357.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 357.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 357.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 357.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 348.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 348.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 347.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 347.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 347.186 38.59 348.334 ;
      VIA 37.776 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 348.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 348.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 347.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 347.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 338.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 337.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 337.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 337.106 38.59 338.254 ;
      VIA 37.776 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 338.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 337.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 337.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 327.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 327.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 327.026 38.59 328.174 ;
      VIA 37.776 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 327.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 327.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 317.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 317.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 316.946 38.59 318.094 ;
      VIA 37.776 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 317.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 317.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 307.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 307.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 306.866 38.59 308.014 ;
      VIA 37.776 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 307.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 307.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 297.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 296.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 296.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 296.786 38.59 297.934 ;
      VIA 37.776 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 297.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 296.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 297.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 287.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 286.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 286.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 286.706 38.59 287.854 ;
      VIA 37.776 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 287.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 286.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 287.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 277.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 276.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 276.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 276.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 276.626 38.59 277.774 ;
      VIA 37.776 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 277.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 276.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 276.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 277.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 267.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 266.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 266.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 266.546 38.59 267.694 ;
      VIA 37.776 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 267.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 266.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 267.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 257.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 256.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 256.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 256.466 38.59 257.614 ;
      VIA 37.776 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 257.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 256.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 257.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 247.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 247.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 247.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 246.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 246.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 246.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 246.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 246.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 246.386 38.59 247.534 ;
      VIA 37.776 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 247.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 247.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 247.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 246.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 246.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 246.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 246.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 246.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 237.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 237.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 237.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 236.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 236.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 236.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 236.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 236.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 236.306 38.59 237.454 ;
      VIA 37.776 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 237.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 237.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 237.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 236.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 236.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 236.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 236.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 236.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 227.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 227.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 226.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 226.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 226.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 226.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 226.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 226.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 226.226 38.59 227.374 ;
      VIA 37.776 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 227.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 227.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 226.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 226.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 226.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 226.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 226.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 226.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 217.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 216.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 216.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 216.146 38.59 217.294 ;
      VIA 37.776 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 217.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 216.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 216.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 207.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 206.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 206.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 206.066 38.59 207.214 ;
      VIA 37.776 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 207.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 206.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 206.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 196.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 196.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 195.986 38.59 197.134 ;
      VIA 37.776 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 196.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 196.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 186.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 186.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 185.906 38.59 187.054 ;
      VIA 37.776 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 186.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 186.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 176.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 176.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 175.826 38.59 176.974 ;
      VIA 37.776 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 176.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 176.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 166.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 165.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 165.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 165.746 38.59 166.894 ;
      VIA 37.776 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 166.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 165.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 166.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 156.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 156.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 156.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 156.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 156.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 155.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 155.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 155.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 155.666 38.59 156.814 ;
      VIA 37.776 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 156.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 156.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 156.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 156.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 156.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 155.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 155.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 156.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 146.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 146.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 146.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 146.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 146.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 145.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 145.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 145.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 145.586 38.59 146.734 ;
      VIA 37.776 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 146.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 146.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 146.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 146.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 146.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 145.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 145.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 146.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 136.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 136.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 136.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 136.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 135.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 135.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 135.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 135.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 135.506 38.59 136.654 ;
      VIA 37.776 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 136.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 136.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 136.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 136.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 135.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 135.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 135.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 136.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 126.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 126.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 126.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 126 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 125.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 125.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 125.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 125.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 125.426 38.59 126.574 ;
      VIA 37.776 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 126.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 126.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 126.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 126 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 125.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 125.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 125.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 126 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 116.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 116.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 116.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 115.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 115.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 115.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 115.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 115.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 115.346 38.59 116.494 ;
      VIA 37.776 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 116.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 116.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 116.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 115.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 115.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 115.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 115.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 115.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 106.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 106.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 105.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 105.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 105.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 105.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 105.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 105.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 105.266 38.59 106.414 ;
      VIA 37.776 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 106.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 106.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 105.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 105.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 105.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 105.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 105.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 105.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 96.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 96.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 95.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 95.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 95.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 95.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 95.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 95.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 95.186 38.59 96.334 ;
      VIA 37.776 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 96.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 96.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 95.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 95.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 95.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 95.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 95.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 95.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 86.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 85.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 85.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 85.106 38.59 86.254 ;
      VIA 37.776 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 86.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 85.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 85.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 75.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 75.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 75.026 38.59 76.174 ;
      VIA 37.776 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 75.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 75.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 65.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 65.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 64.946 38.59 66.094 ;
      VIA 37.776 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 65.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 65.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 55.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 55.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 54.866 38.59 56.014 ;
      VIA 37.776 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 55.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 55.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 45.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 44.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 44.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 44.786 38.59 45.934 ;
      VIA 37.776 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 45.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 44.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 45.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 35.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 34.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 34.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 34.706 38.59 35.854 ;
      VIA 37.776 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 35.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 34.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 35.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 25.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 25.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 25.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 25.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 25.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 24.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 24.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 24.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 24.626 38.59 25.774 ;
      VIA 37.776 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 25.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 25.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 25.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 25.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 25.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 24.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 24.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 25.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 38.056 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 15.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 38.056 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.928 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.8 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.672 14.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 37.544 14.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  36.45 14.546 38.59 15.694 ;
      VIA 37.776 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 15.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.776 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.648 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.392 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.264 14.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 37.52 15.12 via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  567.84 9.506 572.32 605.374 ;
        RECT  523.04 9.506 527.52 605.374 ;
        RECT  478.24 9.506 482.72 605.374 ;
        RECT  433.44 9.506 437.92 605.374 ;
        RECT  388.64 9.506 393.12 605.374 ;
        RECT  343.84 9.506 348.32 605.374 ;
        RECT  299.04 9.506 303.52 605.374 ;
        RECT  254.24 9.506 258.72 605.374 ;
        RECT  209.44 9.506 213.92 605.374 ;
        RECT  164.64 9.506 169.12 605.374 ;
        RECT  119.84 9.506 124.32 605.374 ;
        RECT  75.04 9.506 79.52 605.374 ;
        RECT  30.24 9.506 34.72 605.374 ;
      LAYER Metal1 ;
        RECT  529.2 594.27 609.84 595.17 ;
        RECT  529.2 584.19 609.84 585.09 ;
        RECT  529.2 574.11 609.84 575.01 ;
        RECT  529.2 564.03 609.84 564.93 ;
        RECT  529.2 553.95 609.84 554.85 ;
        RECT  529.2 543.87 609.84 544.77 ;
        RECT  529.2 533.79 609.84 534.69 ;
        RECT  529.2 523.71 609.84 524.61 ;
        RECT  529.2 513.63 609.84 514.53 ;
        RECT  529.2 503.55 609.84 504.45 ;
        RECT  529.2 493.47 609.84 494.37 ;
        RECT  529.2 483.39 609.84 484.29 ;
        RECT  529.2 473.31 609.84 474.21 ;
        RECT  529.2 463.23 609.84 464.13 ;
        RECT  529.2 453.15 609.84 454.05 ;
        RECT  529.2 443.07 609.84 443.97 ;
        RECT  529.2 432.99 609.84 433.89 ;
        RECT  529.2 422.91 609.84 423.81 ;
        RECT  529.2 412.83 609.84 413.73 ;
        RECT  529.2 402.75 609.84 403.65 ;
        RECT  529.2 392.67 609.84 393.57 ;
        RECT  529.2 382.59 609.84 383.49 ;
        RECT  529.2 372.51 609.84 373.41 ;
        RECT  529.2 251.55 609.84 252.45 ;
        RECT  529.2 241.47 609.84 242.37 ;
        RECT  529.2 231.39 609.84 232.29 ;
        RECT  529.2 221.31 609.84 222.21 ;
        RECT  529.2 211.23 609.84 212.13 ;
        RECT  529.2 201.15 609.84 202.05 ;
        RECT  529.2 191.07 609.84 191.97 ;
        RECT  529.2 180.99 609.84 181.89 ;
        RECT  529.2 170.91 609.84 171.81 ;
        RECT  529.2 160.83 609.84 161.73 ;
        RECT  529.2 150.75 609.84 151.65 ;
        RECT  529.2 140.67 609.84 141.57 ;
        RECT  529.2 130.59 609.84 131.49 ;
        RECT  529.2 120.51 609.84 121.41 ;
        RECT  529.2 110.43 609.84 111.33 ;
        RECT  529.2 100.35 609.84 101.25 ;
        RECT  529.2 90.27 609.84 91.17 ;
        RECT  529.2 80.19 609.84 81.09 ;
        RECT  529.2 70.11 609.84 71.01 ;
        RECT  529.2 60.03 609.84 60.93 ;
        RECT  529.2 49.95 609.84 50.85 ;
        RECT  529.2 39.87 609.84 40.77 ;
        RECT  529.2 29.79 609.84 30.69 ;
        RECT  529.2 19.71 609.84 20.61 ;
        RECT  10.08 604.35 609.84 605.25 ;
        RECT  10.08 594.27 92.96 595.17 ;
        RECT  10.08 584.19 92.96 585.09 ;
        RECT  10.08 574.11 92.96 575.01 ;
        RECT  10.08 564.03 92.96 564.93 ;
        RECT  10.08 553.95 92.96 554.85 ;
        RECT  10.08 543.87 92.96 544.77 ;
        RECT  10.08 533.79 92.96 534.69 ;
        RECT  10.08 523.71 92.96 524.61 ;
        RECT  10.08 513.63 92.96 514.53 ;
        RECT  10.08 503.55 92.96 504.45 ;
        RECT  10.08 493.47 92.96 494.37 ;
        RECT  10.08 483.39 92.96 484.29 ;
        RECT  10.08 473.31 92.96 474.21 ;
        RECT  10.08 463.23 92.96 464.13 ;
        RECT  10.08 453.15 92.96 454.05 ;
        RECT  10.08 443.07 92.96 443.97 ;
        RECT  10.08 432.99 92.96 433.89 ;
        RECT  10.08 422.91 92.96 423.81 ;
        RECT  10.08 412.83 92.96 413.73 ;
        RECT  10.08 402.75 92.96 403.65 ;
        RECT  10.08 392.67 92.96 393.57 ;
        RECT  10.08 382.59 92.96 383.49 ;
        RECT  10.08 372.51 92.96 373.41 ;
        RECT  10.08 362.43 609.84 363.33 ;
        RECT  10.08 352.35 609.84 353.25 ;
        RECT  10.08 342.27 609.84 343.17 ;
        RECT  10.08 332.19 609.84 333.09 ;
        RECT  10.08 322.11 609.84 323.01 ;
        RECT  10.08 312.03 609.84 312.93 ;
        RECT  10.08 301.95 609.84 302.85 ;
        RECT  10.08 291.87 609.84 292.77 ;
        RECT  10.08 281.79 609.84 282.69 ;
        RECT  10.08 271.71 609.84 272.61 ;
        RECT  10.08 261.63 609.84 262.53 ;
        RECT  10.08 251.55 92.96 252.45 ;
        RECT  10.08 241.47 92.96 242.37 ;
        RECT  10.08 231.39 92.96 232.29 ;
        RECT  10.08 221.31 92.96 222.21 ;
        RECT  10.08 211.23 92.96 212.13 ;
        RECT  10.08 201.15 92.96 202.05 ;
        RECT  10.08 191.07 92.96 191.97 ;
        RECT  10.08 180.99 92.96 181.89 ;
        RECT  10.08 170.91 92.96 171.81 ;
        RECT  10.08 160.83 92.96 161.73 ;
        RECT  10.08 150.75 92.96 151.65 ;
        RECT  10.08 140.67 92.96 141.57 ;
        RECT  10.08 130.59 92.96 131.49 ;
        RECT  10.08 120.51 92.96 121.41 ;
        RECT  10.08 110.43 92.96 111.33 ;
        RECT  10.08 100.35 92.96 101.25 ;
        RECT  10.08 90.27 92.96 91.17 ;
        RECT  10.08 80.19 92.96 81.09 ;
        RECT  10.08 70.11 92.96 71.01 ;
        RECT  10.08 60.03 92.96 60.93 ;
        RECT  10.08 49.95 92.96 50.85 ;
        RECT  10.08 39.87 92.96 40.77 ;
        RECT  10.08 29.79 92.96 30.69 ;
        RECT  10.08 19.71 92.96 20.61 ;
        RECT  10.08 9.63 609.84 10.53 ;
      VIA 569.956 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 604.226 571.15 605.374 ;
      VIA 570.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 594.146 571.15 595.294 ;
      VIA 570.336 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 584.066 571.15 585.214 ;
      VIA 570.336 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 573.986 571.15 575.134 ;
      VIA 570.336 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 563.906 571.15 565.054 ;
      VIA 570.336 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 553.826 571.15 554.974 ;
      VIA 570.336 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 543.746 571.15 544.894 ;
      VIA 570.336 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 533.666 571.15 534.814 ;
      VIA 570.336 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 523.586 571.15 524.734 ;
      VIA 570.336 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 513.506 571.15 514.654 ;
      VIA 570.336 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 503.426 571.15 504.574 ;
      VIA 570.336 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 493.346 571.15 494.494 ;
      VIA 570.336 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 483.266 571.15 484.414 ;
      VIA 570.336 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 473.186 571.15 474.334 ;
      VIA 570.336 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 463.106 571.15 464.254 ;
      VIA 570.336 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 453.026 571.15 454.174 ;
      VIA 570.336 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 442.946 571.15 444.094 ;
      VIA 570.336 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 432.866 571.15 434.014 ;
      VIA 570.336 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 422.786 571.15 423.934 ;
      VIA 570.336 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 412.706 571.15 413.854 ;
      VIA 570.336 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 402.626 571.15 403.774 ;
      VIA 570.336 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 392.546 571.15 393.694 ;
      VIA 570.336 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 382.466 571.15 383.614 ;
      VIA 570.336 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 372.386 571.15 373.534 ;
      VIA 570.336 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 362.306 571.15 363.454 ;
      VIA 570.336 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 352.226 571.15 353.374 ;
      VIA 570.336 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 342.146 571.15 343.294 ;
      VIA 570.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 332.066 571.15 333.214 ;
      VIA 570.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 321.986 571.15 323.134 ;
      VIA 570.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 311.906 571.15 313.054 ;
      VIA 570.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 301.826 571.15 302.974 ;
      VIA 570.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 291.746 571.15 292.894 ;
      VIA 570.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 281.666 571.15 282.814 ;
      VIA 570.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 271.586 571.15 272.734 ;
      VIA 570.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 261.506 571.15 262.654 ;
      VIA 570.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 251.426 571.15 252.574 ;
      VIA 570.336 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 241.346 571.15 242.494 ;
      VIA 570.336 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 231.266 571.15 232.414 ;
      VIA 570.336 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 221.186 571.15 222.334 ;
      VIA 570.336 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 211.106 571.15 212.254 ;
      VIA 570.336 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 201.026 571.15 202.174 ;
      VIA 570.336 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 190.946 571.15 192.094 ;
      VIA 570.336 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 180.866 571.15 182.014 ;
      VIA 570.336 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 170.786 571.15 171.934 ;
      VIA 570.336 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 160.706 571.15 161.854 ;
      VIA 570.336 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 150.626 571.15 151.774 ;
      VIA 570.336 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 140.546 571.15 141.694 ;
      VIA 570.336 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 130.466 571.15 131.614 ;
      VIA 570.336 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 120.386 571.15 121.534 ;
      VIA 570.336 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 110.306 571.15 111.454 ;
      VIA 570.336 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 100.226 571.15 101.374 ;
      VIA 570.336 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 90.146 571.15 91.294 ;
      VIA 570.336 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 80.066 571.15 81.214 ;
      VIA 570.336 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 69.986 571.15 71.134 ;
      VIA 570.336 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 59.906 571.15 61.054 ;
      VIA 570.336 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 49.826 571.15 50.974 ;
      VIA 570.336 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 39.746 571.15 40.894 ;
      VIA 570.336 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 29.666 571.15 30.814 ;
      VIA 570.336 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 19.586 571.15 20.734 ;
      VIA 570.336 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 569.956 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.956 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.828 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.7 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.572 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 569.444 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  569.01 9.506 571.15 10.654 ;
      VIA 570.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 569.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 570.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 604.226 526.35 605.374 ;
      VIA 525.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 362.306 526.35 363.454 ;
      VIA 525.536 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 352.226 526.35 353.374 ;
      VIA 525.536 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 342.146 526.35 343.294 ;
      VIA 525.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 332.066 526.35 333.214 ;
      VIA 525.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 321.986 526.35 323.134 ;
      VIA 525.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 311.906 526.35 313.054 ;
      VIA 525.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 301.826 526.35 302.974 ;
      VIA 525.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 291.746 526.35 292.894 ;
      VIA 525.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 281.666 526.35 282.814 ;
      VIA 525.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 271.586 526.35 272.734 ;
      VIA 525.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 261.506 526.35 262.654 ;
      VIA 525.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 525.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 525.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  524.21 9.506 526.35 10.654 ;
      VIA 525.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 525.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 604.226 481.55 605.374 ;
      VIA 480.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 362.306 481.55 363.454 ;
      VIA 480.736 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 352.226 481.55 353.374 ;
      VIA 480.736 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 342.146 481.55 343.294 ;
      VIA 480.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 332.066 481.55 333.214 ;
      VIA 480.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 321.986 481.55 323.134 ;
      VIA 480.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 311.906 481.55 313.054 ;
      VIA 480.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 301.826 481.55 302.974 ;
      VIA 480.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 291.746 481.55 292.894 ;
      VIA 480.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 281.666 481.55 282.814 ;
      VIA 480.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 271.586 481.55 272.734 ;
      VIA 480.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 261.506 481.55 262.654 ;
      VIA 480.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 480.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 480.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  479.41 9.506 481.55 10.654 ;
      VIA 480.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 480.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 604.226 436.75 605.374 ;
      VIA 435.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 362.306 436.75 363.454 ;
      VIA 435.936 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 352.226 436.75 353.374 ;
      VIA 435.936 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 342.146 436.75 343.294 ;
      VIA 435.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 332.066 436.75 333.214 ;
      VIA 435.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 321.986 436.75 323.134 ;
      VIA 435.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 311.906 436.75 313.054 ;
      VIA 435.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 301.826 436.75 302.974 ;
      VIA 435.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 291.746 436.75 292.894 ;
      VIA 435.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 281.666 436.75 282.814 ;
      VIA 435.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 271.586 436.75 272.734 ;
      VIA 435.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 261.506 436.75 262.654 ;
      VIA 435.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 435.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 435.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  434.61 9.506 436.75 10.654 ;
      VIA 435.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 435.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 604.226 391.95 605.374 ;
      VIA 391.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 362.306 391.95 363.454 ;
      VIA 391.136 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 352.226 391.95 353.374 ;
      VIA 391.136 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 342.146 391.95 343.294 ;
      VIA 391.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 332.066 391.95 333.214 ;
      VIA 391.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 321.986 391.95 323.134 ;
      VIA 391.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 311.906 391.95 313.054 ;
      VIA 391.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 301.826 391.95 302.974 ;
      VIA 391.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 291.746 391.95 292.894 ;
      VIA 391.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 281.666 391.95 282.814 ;
      VIA 391.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 271.586 391.95 272.734 ;
      VIA 391.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 261.506 391.95 262.654 ;
      VIA 391.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 390.856 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.856 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.728 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.6 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.472 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 390.344 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  389.81 9.506 391.95 10.654 ;
      VIA 391.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 391.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 390.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 604.226 347.15 605.374 ;
      VIA 346.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 362.306 347.15 363.454 ;
      VIA 346.336 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 352.226 347.15 353.374 ;
      VIA 346.336 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 342.146 347.15 343.294 ;
      VIA 346.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 332.066 347.15 333.214 ;
      VIA 346.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 321.986 347.15 323.134 ;
      VIA 346.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 311.906 347.15 313.054 ;
      VIA 346.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 301.826 347.15 302.974 ;
      VIA 346.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 291.746 347.15 292.894 ;
      VIA 346.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 281.666 347.15 282.814 ;
      VIA 346.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 271.586 347.15 272.734 ;
      VIA 346.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 261.506 347.15 262.654 ;
      VIA 346.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 346.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 346.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  345.01 9.506 347.15 10.654 ;
      VIA 346.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 345.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 346.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 604.226 302.35 605.374 ;
      VIA 301.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 362.306 302.35 363.454 ;
      VIA 301.536 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 352.226 302.35 353.374 ;
      VIA 301.536 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 342.146 302.35 343.294 ;
      VIA 301.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 332.066 302.35 333.214 ;
      VIA 301.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 321.986 302.35 323.134 ;
      VIA 301.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 311.906 302.35 313.054 ;
      VIA 301.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 301.826 302.35 302.974 ;
      VIA 301.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 291.746 302.35 292.894 ;
      VIA 301.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 281.666 302.35 282.814 ;
      VIA 301.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 271.586 302.35 272.734 ;
      VIA 301.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 261.506 302.35 262.654 ;
      VIA 301.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 301.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 301.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  300.21 9.506 302.35 10.654 ;
      VIA 301.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 301.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 604.226 257.55 605.374 ;
      VIA 256.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 362.306 257.55 363.454 ;
      VIA 256.736 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 352.226 257.55 353.374 ;
      VIA 256.736 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 342.146 257.55 343.294 ;
      VIA 256.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 332.066 257.55 333.214 ;
      VIA 256.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 321.986 257.55 323.134 ;
      VIA 256.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 311.906 257.55 313.054 ;
      VIA 256.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 301.826 257.55 302.974 ;
      VIA 256.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 291.746 257.55 292.894 ;
      VIA 256.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 281.666 257.55 282.814 ;
      VIA 256.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 271.586 257.55 272.734 ;
      VIA 256.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 261.506 257.55 262.654 ;
      VIA 256.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 256.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 256.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  255.41 9.506 257.55 10.654 ;
      VIA 256.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 256.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 604.226 212.75 605.374 ;
      VIA 211.936 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 362.306 212.75 363.454 ;
      VIA 211.936 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 352.226 212.75 353.374 ;
      VIA 211.936 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 342.146 212.75 343.294 ;
      VIA 211.936 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 332.066 212.75 333.214 ;
      VIA 211.936 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 321.986 212.75 323.134 ;
      VIA 211.936 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 311.906 212.75 313.054 ;
      VIA 211.936 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 301.826 212.75 302.974 ;
      VIA 211.936 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 291.746 212.75 292.894 ;
      VIA 211.936 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 281.666 212.75 282.814 ;
      VIA 211.936 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 271.586 212.75 272.734 ;
      VIA 211.936 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 261.506 212.75 262.654 ;
      VIA 211.936 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 211.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 211.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  210.61 9.506 212.75 10.654 ;
      VIA 211.936 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.936 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.808 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.552 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.424 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 211.68 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 604.226 167.95 605.374 ;
      VIA 167.136 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 362.306 167.95 363.454 ;
      VIA 167.136 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 352.226 167.95 353.374 ;
      VIA 167.136 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 342.146 167.95 343.294 ;
      VIA 167.136 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 332.066 167.95 333.214 ;
      VIA 167.136 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 321.986 167.95 323.134 ;
      VIA 167.136 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 311.906 167.95 313.054 ;
      VIA 167.136 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 301.826 167.95 302.974 ;
      VIA 167.136 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 291.746 167.95 292.894 ;
      VIA 167.136 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 281.666 167.95 282.814 ;
      VIA 167.136 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 271.586 167.95 272.734 ;
      VIA 167.136 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 261.506 167.95 262.654 ;
      VIA 167.136 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 166.756 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.756 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.628 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.5 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.372 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 166.244 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  165.81 9.506 167.95 10.654 ;
      VIA 167.136 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.136 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 167.008 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.752 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.624 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 166.88 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 604.226 123.15 605.374 ;
      VIA 122.336 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 362.306 123.15 363.454 ;
      VIA 122.336 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 352.226 123.15 353.374 ;
      VIA 122.336 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 342.146 123.15 343.294 ;
      VIA 122.336 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 332.066 123.15 333.214 ;
      VIA 122.336 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 321.986 123.15 323.134 ;
      VIA 122.336 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 311.906 123.15 313.054 ;
      VIA 122.336 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 301.826 123.15 302.974 ;
      VIA 122.336 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 291.746 123.15 292.894 ;
      VIA 122.336 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 281.666 123.15 282.814 ;
      VIA 122.336 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 271.586 123.15 272.734 ;
      VIA 122.336 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 261.506 123.15 262.654 ;
      VIA 122.336 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 122.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 122.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  121.01 9.506 123.15 10.654 ;
      VIA 122.336 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.336 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.208 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.952 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 121.824 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 122.08 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 604.226 78.35 605.374 ;
      VIA 77.536 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 594.146 78.35 595.294 ;
      VIA 77.536 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 584.066 78.35 585.214 ;
      VIA 77.536 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 573.986 78.35 575.134 ;
      VIA 77.536 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 563.906 78.35 565.054 ;
      VIA 77.536 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 553.826 78.35 554.974 ;
      VIA 77.536 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 543.746 78.35 544.894 ;
      VIA 77.536 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 533.666 78.35 534.814 ;
      VIA 77.536 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 523.586 78.35 524.734 ;
      VIA 77.536 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 513.506 78.35 514.654 ;
      VIA 77.536 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 503.426 78.35 504.574 ;
      VIA 77.536 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 493.346 78.35 494.494 ;
      VIA 77.536 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 483.266 78.35 484.414 ;
      VIA 77.536 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 473.186 78.35 474.334 ;
      VIA 77.536 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 463.106 78.35 464.254 ;
      VIA 77.536 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 453.026 78.35 454.174 ;
      VIA 77.536 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 442.946 78.35 444.094 ;
      VIA 77.536 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 432.866 78.35 434.014 ;
      VIA 77.536 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 422.786 78.35 423.934 ;
      VIA 77.536 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 412.706 78.35 413.854 ;
      VIA 77.536 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 402.626 78.35 403.774 ;
      VIA 77.536 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 392.546 78.35 393.694 ;
      VIA 77.536 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 382.466 78.35 383.614 ;
      VIA 77.536 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 372.386 78.35 373.534 ;
      VIA 77.536 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 362.306 78.35 363.454 ;
      VIA 77.536 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 352.226 78.35 353.374 ;
      VIA 77.536 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 342.146 78.35 343.294 ;
      VIA 77.536 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 332.066 78.35 333.214 ;
      VIA 77.536 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 321.986 78.35 323.134 ;
      VIA 77.536 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 311.906 78.35 313.054 ;
      VIA 77.536 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 301.826 78.35 302.974 ;
      VIA 77.536 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 291.746 78.35 292.894 ;
      VIA 77.536 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 281.666 78.35 282.814 ;
      VIA 77.536 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 271.586 78.35 272.734 ;
      VIA 77.536 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 261.506 78.35 262.654 ;
      VIA 77.536 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 251.426 78.35 252.574 ;
      VIA 77.536 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 241.346 78.35 242.494 ;
      VIA 77.536 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 231.266 78.35 232.414 ;
      VIA 77.536 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 221.186 78.35 222.334 ;
      VIA 77.536 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 211.106 78.35 212.254 ;
      VIA 77.536 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 201.026 78.35 202.174 ;
      VIA 77.536 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 190.946 78.35 192.094 ;
      VIA 77.536 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 180.866 78.35 182.014 ;
      VIA 77.536 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 170.786 78.35 171.934 ;
      VIA 77.536 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 160.706 78.35 161.854 ;
      VIA 77.536 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 150.626 78.35 151.774 ;
      VIA 77.536 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 140.546 78.35 141.694 ;
      VIA 77.536 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 130.466 78.35 131.614 ;
      VIA 77.536 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 120.386 78.35 121.534 ;
      VIA 77.536 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 110.306 78.35 111.454 ;
      VIA 77.536 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 100.226 78.35 101.374 ;
      VIA 77.536 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 90.146 78.35 91.294 ;
      VIA 77.536 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 80.066 78.35 81.214 ;
      VIA 77.536 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 69.986 78.35 71.134 ;
      VIA 77.536 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 59.906 78.35 61.054 ;
      VIA 77.536 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 49.826 78.35 50.974 ;
      VIA 77.536 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 39.746 78.35 40.894 ;
      VIA 77.536 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 29.666 78.35 30.814 ;
      VIA 77.536 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 19.586 78.35 20.734 ;
      VIA 77.536 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 77.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 77.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  76.21 9.506 78.35 10.654 ;
      VIA 77.536 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.536 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.408 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.152 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.024 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 77.28 10.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 605.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 605.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 604.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 604.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 604.226 33.55 605.374 ;
      VIA 32.736 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 605.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 605.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 604.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 604.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 595.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 594.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 594.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 594.146 33.55 595.294 ;
      VIA 32.736 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 595.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 594.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 594.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 585.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 584.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 584.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 584.066 33.55 585.214 ;
      VIA 32.736 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 585.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 584.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 584.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 574.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 574.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 573.986 33.55 575.134 ;
      VIA 32.736 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 574.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 574.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 564.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 564.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 563.906 33.55 565.054 ;
      VIA 32.736 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 564.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 564.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 554.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 554.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 553.826 33.55 554.974 ;
      VIA 32.736 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 554.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 554.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 544.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 543.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 543.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 543.746 33.55 544.894 ;
      VIA 32.736 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 544.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 543.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 544.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 534.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 534.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 534.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 534.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 534.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 533.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 533.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 533.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 533.666 33.55 534.814 ;
      VIA 32.736 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 534.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 534.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 534.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 534.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 534.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 533.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 533.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 534.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 524.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 524.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 524.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 524.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 524.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 523.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 523.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 523.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 523.586 33.55 524.734 ;
      VIA 32.736 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 524.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 524.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 524.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 524.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 524.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 523.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 523.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 524.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 514.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 514.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 514.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 514.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 513.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 513.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 513.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 513.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 513.506 33.55 514.654 ;
      VIA 32.736 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 514.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 514.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 514.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 514.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 513.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 513.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 513.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 514.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 504.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 504.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 504.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 503.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 503.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 503.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 503.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 503.426 33.55 504.574 ;
      VIA 32.736 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 504.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 504.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 504.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 503.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 503.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 503.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 504 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 494.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 494.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 494.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 493.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 493.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 493.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 493.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 493.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 493.346 33.55 494.494 ;
      VIA 32.736 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 494.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 494.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 494.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 493.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 493.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 493.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 493.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 493.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 484.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 484.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 483.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 483.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 483.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 483.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 483.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 483.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 483.266 33.55 484.414 ;
      VIA 32.736 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 484.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 484.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 483.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 483.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 483.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 483.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 483.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 483.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 474.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 474.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 473.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 473.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 473.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 473.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 473.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 473.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 473.186 33.55 474.334 ;
      VIA 32.736 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 474.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 474.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 473.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 473.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 473.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 473.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 473.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 473.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 464.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 463.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 463.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 463.106 33.55 464.254 ;
      VIA 32.736 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 464.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 463.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 463.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 453.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 453.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 453.026 33.55 454.174 ;
      VIA 32.736 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 453.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 453.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 443.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 443.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 442.946 33.55 444.094 ;
      VIA 32.736 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 443.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 443.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 433.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 433.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 432.866 33.55 434.014 ;
      VIA 32.736 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 433.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 433.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 423.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 422.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 422.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 422.786 33.55 423.934 ;
      VIA 32.736 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 423.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 422.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 423.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 413.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 412.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 412.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 412.706 33.55 413.854 ;
      VIA 32.736 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 413.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 412.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 413.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 403.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 403.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 403.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 403.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 403.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 402.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 402.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 402.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 402.626 33.55 403.774 ;
      VIA 32.736 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 403.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 403.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 403.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 403.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 403.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 402.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 402.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 403.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 393.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 393.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 393.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 393.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 392.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 392.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 392.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 392.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 392.546 33.55 393.694 ;
      VIA 32.736 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 393.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 393.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 393.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 393.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 392.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 392.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 392.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 393.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 383.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 383.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 383.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 383.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 382.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 382.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 382.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 382.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 382.466 33.55 383.614 ;
      VIA 32.736 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 383.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 383.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 383.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 383.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 382.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 382.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 382.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 383.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 373.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 373.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 373.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 372.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 372.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 372.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 372.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 372.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 372.386 33.55 373.534 ;
      VIA 32.736 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 373.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 373.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 373.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 372.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 372.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 372.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 372.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 372.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 363.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 363.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 363.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 362.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 362.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 362.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 362.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 362.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 362.306 33.55 363.454 ;
      VIA 32.736 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 363.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 363.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 363.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 362.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 362.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 362.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 362.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 362.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 353.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 353.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 352.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 352.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 352.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 352.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 352.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 352.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 352.226 33.55 353.374 ;
      VIA 32.736 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 353.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 353.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 352.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 352.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 352.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 352.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 352.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 352.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 343.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 342.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 342.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 342.146 33.55 343.294 ;
      VIA 32.736 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 343.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 342.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 342.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 333.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 332.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 332.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 332.066 33.55 333.214 ;
      VIA 32.736 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 333.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 332.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 332.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 322.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 322.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 321.986 33.55 323.134 ;
      VIA 32.736 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 322.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 322.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 312.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 312.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 311.906 33.55 313.054 ;
      VIA 32.736 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 312.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 312.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 302.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 302.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 301.826 33.55 302.974 ;
      VIA 32.736 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 302.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 302.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 292.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 291.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 291.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 291.746 33.55 292.894 ;
      VIA 32.736 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 292.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 291.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 292.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 282.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 281.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 281.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 281.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 281.666 33.55 282.814 ;
      VIA 32.736 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 282.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 281.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 281.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 282.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 272.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 271.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 271.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 271.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 271.586 33.55 272.734 ;
      VIA 32.736 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 272.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 271.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 271.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 272.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 262.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 261.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 261.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 261.506 33.55 262.654 ;
      VIA 32.736 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 262.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 261.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 262.08 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 252.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 252.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 252.128 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 252 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 251.872 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 251.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 251.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 251.616 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 251.426 33.55 252.574 ;
      VIA 32.736 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 252.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 252.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 252.128 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 252 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 251.872 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 251.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 251.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 252 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 242.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 242.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 242.048 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 241.92 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 241.792 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 241.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 241.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 241.536 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 241.346 33.55 242.494 ;
      VIA 32.736 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 242.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 242.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 242.048 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 241.92 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 241.792 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 241.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 241.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 241.92 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 232.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 232.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 231.968 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 231.84 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 231.712 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 231.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 231.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 231.456 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 231.266 33.55 232.414 ;
      VIA 32.736 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 232.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 232.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 231.968 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 231.84 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 231.712 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 231.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 231.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 231.84 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 222.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 222.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 221.888 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 221.76 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 221.632 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 221.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 221.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 221.376 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 221.186 33.55 222.334 ;
      VIA 32.736 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 222.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 222.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 221.888 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 221.76 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 221.632 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 221.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 221.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 221.76 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 212.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.808 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.68 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.552 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 211.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 211.296 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 211.106 33.55 212.254 ;
      VIA 32.736 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 212.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.808 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.68 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.552 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 211.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 211.68 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.728 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.6 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.472 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 201.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 201.216 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 201.026 33.55 202.174 ;
      VIA 32.736 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.728 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.6 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.472 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 201.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 201.6 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.648 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.52 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.392 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 191.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 191.136 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 190.946 33.55 192.094 ;
      VIA 32.736 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.648 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.52 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.392 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 191.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 191.52 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.568 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.44 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.312 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 181.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 181.056 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 180.866 33.55 182.014 ;
      VIA 32.736 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.568 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.44 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.312 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 181.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 181.44 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.744 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.616 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.488 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.36 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.232 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 171.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 170.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 170.976 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 170.786 33.55 171.934 ;
      VIA 32.736 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.744 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.616 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.488 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.36 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.232 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 171.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 170.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 171.36 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.664 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.536 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.408 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.28 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.152 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 161.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 160.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 160.896 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 160.706 33.55 161.854 ;
      VIA 32.736 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.664 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.536 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.408 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.28 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.152 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 161.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 160.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 161.28 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 151.584 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 151.456 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 151.328 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 151.2 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 151.072 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 150.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 150.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 150.816 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 150.626 33.55 151.774 ;
      VIA 32.736 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 151.584 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 151.456 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 151.328 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 151.2 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 151.072 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 150.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 150.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 151.2 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 141.504 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 141.376 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 141.248 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 141.12 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 140.992 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 140.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 140.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 140.736 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 140.546 33.55 141.694 ;
      VIA 32.736 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 141.504 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 141.376 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 141.248 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 141.12 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 140.992 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 140.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 140.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 141.12 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 131.424 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 131.296 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 131.168 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 131.04 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 130.912 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 130.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 130.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 130.656 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 130.466 33.55 131.614 ;
      VIA 32.736 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 131.424 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 131.296 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 131.168 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 131.04 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 130.912 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 130.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 130.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 131.04 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 121.344 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 121.216 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 121.088 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 120.96 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 120.832 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 120.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 120.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 120.576 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 120.386 33.55 121.534 ;
      VIA 32.736 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 121.344 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 121.216 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 121.088 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 120.96 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 120.832 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 120.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 120.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 120.96 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 111.264 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 111.136 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 111.008 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 110.88 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 110.752 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 110.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 110.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 110.496 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 110.306 33.55 111.454 ;
      VIA 32.736 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 111.264 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 111.136 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 111.008 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 110.88 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 110.752 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 110.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 110.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 110.88 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 101.184 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 101.056 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 100.928 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 100.8 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 100.672 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 100.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 100.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 100.416 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 100.226 33.55 101.374 ;
      VIA 32.736 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 101.184 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 101.056 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 100.928 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 100.8 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 100.672 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 100.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 100.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 100.8 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 91.104 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.976 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.848 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.72 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.592 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 90.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 90.336 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 90.146 33.55 91.294 ;
      VIA 32.736 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 91.104 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.976 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.848 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.72 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.592 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 90.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 90.72 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 81.024 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.896 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.768 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.64 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.512 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.384 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 80.256 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 80.256 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 80.066 33.55 81.214 ;
      VIA 32.736 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 81.024 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.896 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.768 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.64 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.512 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.384 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 80.256 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 80.64 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.944 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.816 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.688 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.56 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.432 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.304 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 70.176 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 70.176 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 69.986 33.55 71.134 ;
      VIA 32.736 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.944 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.816 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.688 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.56 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.432 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.304 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 70.176 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 70.56 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.864 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.736 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.608 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.48 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.352 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.224 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 60.096 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 60.096 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 59.906 33.55 61.054 ;
      VIA 32.736 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.864 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.736 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.608 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.48 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.352 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.224 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 60.096 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 60.48 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.784 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.656 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.528 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.4 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.272 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.144 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 50.016 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 50.016 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 49.826 33.55 50.974 ;
      VIA 32.736 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.784 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.656 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.528 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.4 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.272 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.144 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 50.016 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 50.4 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.704 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.576 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.448 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.32 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.192 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 40.064 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 39.936 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 39.936 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 39.746 33.55 40.894 ;
      VIA 32.736 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.704 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.576 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.448 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.32 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.192 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 40.064 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 39.936 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 40.32 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 30.624 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 30.496 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 30.368 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 30.24 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 30.112 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 29.984 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 29.856 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 29.856 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 29.666 33.55 30.814 ;
      VIA 32.736 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 30.624 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 30.496 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 30.368 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 30.24 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 30.112 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 29.984 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 29.856 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 30.24 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 20.544 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 20.416 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 20.288 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 20.16 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 20.032 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 19.904 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 19.776 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 19.776 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 19.586 33.55 20.734 ;
      VIA 32.736 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 20.544 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 20.416 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 20.288 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 20.16 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 20.032 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 19.904 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 19.776 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 20.16 via1_2_8960_1800_1_4_1240_1240 ;
      VIA 32.656 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.464 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.336 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.208 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 10.08 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.952 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.824 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.656 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.528 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.4 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.272 9.696 via3_4_8960_1800_1_1_256_256 ;
      VIA 32.144 9.696 via3_4_8960_1800_1_1_256_256 ;
      LAYER Metal2 ;
        RECT  31.41 9.506 33.55 10.654 ;
      VIA 32.736 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.464 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.336 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.208 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 10.08 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.952 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.824 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.736 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.608 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.352 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.224 9.696 via2_3_8960_1800_1_1_256_256 ;
      VIA 32.48 10.08 via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VSS
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  267.08 0 267.52 1.28 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  258.08 0 258.52 1.28 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  249.08 0 249.52 1.28 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  376.88 0 377.32 1.28 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  371.48 0 371.92 1.28 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  367.88 0 368.32 1.28 ;
    END
  END addr[5]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  360.68 0 361.12 1.28 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  234.68 0 235.12 1.28 ;
    END
  END clk
  PIN idat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  105.08 0 105.52 1.28 ;
    END
  END idat[0]
  PIN idat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 364.42 0.52 364.7 ;
    END
  END idat[10]
  PIN idat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 368.9 0.52 369.18 ;
    END
  END idat[11]
  PIN idat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 364.42 620 364.7 ;
    END
  END idat[12]
  PIN idat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 368.9 620 369.18 ;
    END
  END idat[13]
  PIN idat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 371.14 620 371.42 ;
    END
  END idat[14]
  PIN idat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 366.66 620 366.94 ;
    END
  END idat[15]
  PIN idat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  155.48 0 155.92 1.28 ;
    END
  END idat[1]
  PIN idat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  162.68 0 163.12 1.28 ;
    END
  END idat[2]
  PIN idat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  214.88 0 215.32 1.28 ;
    END
  END idat[3]
  PIN idat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  402.08 0 402.52 1.28 ;
    END
  END idat[4]
  PIN idat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  454.28 0 454.72 1.28 ;
    END
  END idat[5]
  PIN idat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  459.68 0 460.12 1.28 ;
    END
  END idat[6]
  PIN idat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  511.88 0 512.32 1.28 ;
    END
  END idat[7]
  PIN idat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 370.02 0.52 370.3 ;
    END
  END idat[8]
  PIN idat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 367.78 0.52 368.06 ;
    END
  END idat[9]
  PIN odat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  112.28 0 112.72 1.28 ;
    END
  END odat[0]
  PIN odat[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 371.14 0.52 371.42 ;
    END
  END odat[10]
  PIN odat[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 372.26 0.52 372.54 ;
    END
  END odat[11]
  PIN odat[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 365.54 620 365.82 ;
    END
  END odat[12]
  PIN odat[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 370.02 620 370.3 ;
    END
  END odat[13]
  PIN odat[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 372.26 620 372.54 ;
    END
  END odat[14]
  PIN odat[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  619.48 367.78 620 368.06 ;
    END
  END odat[15]
  PIN odat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  153.68 0 154.12 1.28 ;
    END
  END odat[1]
  PIN odat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  166.28 0 166.72 1.28 ;
    END
  END odat[2]
  PIN odat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  205.88 0 206.32 1.28 ;
    END
  END odat[3]
  PIN odat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  409.28 0 409.72 1.28 ;
    END
  END odat[4]
  PIN odat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  450.68 0 451.12 1.28 ;
    END
  END odat[5]
  PIN odat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  463.28 0 463.72 1.28 ;
    END
  END odat[6]
  PIN odat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  504.68 0 505.12 1.28 ;
    END
  END odat[7]
  PIN odat[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 365.54 0.52 365.82 ;
    END
  END odat[8]
  PIN odat[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT  0 366.66 0.52 366.94 ;
    END
  END odat[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  297.68 0 298.12 1.28 ;
    END
  END we
  OBS
    LAYER Metal1 ;
     RECT  10.08 9.63 93.965 610.29 ;
     RECT  93.965 8.845 112.445 610.29 ;
     RECT  112.445 8.285 117.715 610.29 ;
     RECT  117.715 8.845 159.485 610.29 ;
     RECT  159.485 8.285 272.835 610.29 ;
     RECT  272.835 8.845 277.875 610.29 ;
     RECT  277.875 9.63 304.525 610.29 ;
     RECT  304.525 8.845 350.675 610.29 ;
     RECT  350.675 9.63 371.165 610.29 ;
     RECT  371.165 8.285 408.685 610.29 ;
     RECT  408.685 7.725 409.245 610.29 ;
     RECT  409.245 7.165 419.555 610.29 ;
     RECT  419.555 8.285 460.205 610.29 ;
     RECT  460.205 7.725 476.675 610.29 ;
     RECT  476.675 8.285 532.675 610.29 ;
     RECT  532.675 8.845 533.795 610.29 ;
     RECT  533.795 9.63 609.84 610.29 ;
    LAYER Metal2 ;
     RECT  112.42 8.07 112.7 8.26 ;
     RECT  460.18 7.7 460.46 8.26 ;
     RECT  418.18 8.26 420.14 8.54 ;
     RECT  259.14 8.26 272.86 8.63 ;
     RECT  383.46 8.26 383.74 8.63 ;
     RECT  167.86 8.26 168.14 8.82 ;
     RECT  251.86 8.63 272.86 8.82 ;
     RECT  377.86 8.63 383.74 8.82 ;
     RECT  532.42 8.26 532.7 8.82 ;
     RECT  93.94 8.82 94.22 9.38 ;
     RECT  112.42 8.26 117.74 9.38 ;
     RECT  167.86 8.82 173.18 9.38 ;
     RECT  205.94 6.58 206.22 9.38 ;
     RECT  304.5 8.82 304.78 9.38 ;
     RECT  350.42 8.82 392.7 9.38 ;
     RECT  409.78 8.63 417.9 9.38 ;
     RECT  456.82 8.26 460.46 9.38 ;
     RECT  93.94 9.38 117.74 9.506 ;
     RECT  350.42 9.38 417.9 9.506 ;
     RECT  476.42 7.7 476.7 9.506 ;
     RECT  532.42 8.82 533.82 9.506 ;
     RECT  157.5 9.38 173.18 11.34 ;
     RECT  434.61 9.506 436.75 11.34 ;
     RECT  456.82 9.38 461.3 11.34 ;
     RECT  157.5 11.34 180.685 11.62 ;
     RECT  434.61 11.34 461.3 11.62 ;
     RECT  476.42 9.506 481.55 11.62 ;
     RECT  524.21 9.506 533.82 11.62 ;
     RECT  205.94 9.38 216.02 12.18 ;
     RECT  147.98 11.62 180.685 12.31 ;
     RECT  506.445 11.34 506.725 12.31 ;
     RECT  520.66 11.62 533.82 12.31 ;
     RECT  236.18 12.46 236.46 12.74 ;
     RECT  251.86 8.82 277.9 12.74 ;
     RECT  434.61 11.62 481.55 12.74 ;
     RECT  200.62 12.18 216.02 13.02 ;
     RECT  93.94 9.506 123.15 13.3 ;
     RECT  506.445 12.31 533.82 13.3 ;
     RECT  31.41 9.506 33.55 14.546 ;
     RECT  76.21 9.506 78.35 14.546 ;
     RECT  90.02 13.3 123.15 14.546 ;
     RECT  138.46 12.31 180.685 14.546 ;
     RECT  298.62 9.38 304.78 14.546 ;
     RECT  434.61 12.74 485.94 14.546 ;
     RECT  569.01 9.506 571.15 14.546 ;
     RECT  236.18 12.74 282.1 16.66 ;
     RECT  506.445 13.3 537.74 16.66 ;
     RECT  76.21 14.546 180.685 20 ;
     RECT  200.62 13.02 221.9 20 ;
     RECT  235.06 16.66 282.1 20 ;
     RECT  298.62 14.546 307.39 20 ;
     RECT  345.01 9.506 417.9 20 ;
     RECT  434.61 14.546 486.59 20 ;
     RECT  504.98 16.66 537.74 20 ;
     RECT  76.21 20 537.74 252.88 ;
     RECT  236.18 252.88 262.59 259.98 ;
     RECT  117.46 252.88 128.19 260.4 ;
     RECT  208.74 252.88 217.79 263.34 ;
     RECT  236.18 259.98 243.74 263.34 ;
     RECT  236.18 263.34 236.46 274.82 ;
     RECT  255.41 259.98 262.59 274.82 ;
     RECT  242.9 274.82 262.59 275.1 ;
     RECT  210.61 263.34 217.79 348.74 ;
     RECT  255.41 275.1 262.59 348.74 ;
     RECT  300.21 252.88 307.39 348.74 ;
     RECT  76.21 252.88 94.22 349.02 ;
     RECT  76.21 349.02 90.86 349.58 ;
     RECT  76.21 349.58 88.06 350.42 ;
     RECT  165.81 252.88 172.99 350.42 ;
     RECT  367.78 349.3 368.06 350.42 ;
     RECT  208.74 348.74 217.79 350.79 ;
     RECT  242.9 275.1 243.18 350.79 ;
     RECT  207.62 350.79 217.79 350.98 ;
     RECT  367.78 350.42 371.42 350.98 ;
     RECT  434.61 252.88 441.79 350.98 ;
     RECT  235.06 350.79 243.18 351.12 ;
     RECT  156.1 350.42 172.99 351.54 ;
     RECT  242.9 351.12 243.18 351.54 ;
     RECT  255.41 348.74 266.7 351.54 ;
     RECT  410.9 348.74 411.74 351.54 ;
     RECT  464.1 350.42 464.38 353.59 ;
     RECT  479.41 252.88 486.59 353.59 ;
     RECT  434.61 350.98 451.5 353.78 ;
     RECT  464.1 353.59 486.59 353.78 ;
     RECT  599.06 351.54 599.34 354.34 ;
     RECT  524.21 252.88 537.74 354.9 ;
     RECT  596.82 354.34 599.34 354.9 ;
     RECT  13.86 351.54 14.14 355.46 ;
     RECT  31.41 14.546 38.59 355.46 ;
     RECT  389.81 252.88 396.99 355.46 ;
     RECT  410.34 351.54 411.74 355.46 ;
     RECT  512.82 354.9 537.74 355.46 ;
     RECT  569.01 14.546 576.19 355.46 ;
     RECT  109.06 355.46 109.34 355.83 ;
     RECT  121.01 260.4 128.19 355.83 ;
     RECT  596.82 354.9 604.38 356.02 ;
     RECT  434.61 353.78 486.59 356.16 ;
     RECT  504.98 355.46 537.74 356.39 ;
     RECT  596.82 356.02 604.94 356.58 ;
     RECT  58.66 356.39 58.94 356.72 ;
     RECT  499.38 356.39 537.74 356.72 ;
     RECT  109.06 355.83 128.19 359.94 ;
     RECT  13.86 355.46 38.59 360.78 ;
     RECT  13.02 360.78 38.59 361.06 ;
     RECT  389.81 355.46 411.74 361.34 ;
     RECT  596.82 356.58 606.06 363.3 ;
     RECT  242.9 351.54 266.7 364.98 ;
     RECT  70.98 350.42 88.06 366.1 ;
     RECT  70.98 366.1 93.66 367.22 ;
     RECT  108.5 359.94 128.19 367.22 ;
     RECT  70.98 367.22 128.19 368 ;
     RECT  152.74 351.54 172.99 368 ;
     RECT  206.5 350.98 217.79 368 ;
     RECT  235.34 364.98 266.7 368 ;
     RECT  298.34 348.74 307.39 368 ;
     RECT  345.01 252.88 352.19 368 ;
     RECT  367.78 350.98 377.02 368 ;
     RECT  389.81 361.34 412.525 368 ;
     RECT  434.61 356.16 464.38 368 ;
     RECT  479.41 356.16 486.59 368 ;
     RECT  504.98 356.72 537.74 368 ;
     RECT  596.82 363.3 615.58 368.62 ;
     RECT  596.82 368.62 606.06 369.46 ;
     RECT  70.98 368 537.74 370.3 ;
     RECT  569.01 355.46 579.74 370.58 ;
     RECT  596.26 369.46 606.06 370.58 ;
     RECT  569.01 370.58 606.06 370.86 ;
     RECT  590.38 370.86 606.06 375.06 ;
     RECT  596.26 375.06 606.06 376.18 ;
     RECT  12.18 361.06 38.59 377.58 ;
     RECT  598.5 376.18 606.06 380.1 ;
     RECT  76.21 370.3 537.74 380.38 ;
     RECT  95 380.38 537.74 380.94 ;
     RECT  13.02 377.58 38.59 382.62 ;
     RECT  13.02 382.62 18.9 385.14 ;
     RECT  95 380.94 537.18 385.42 ;
     RECT  598.5 380.1 605.78 385.42 ;
     RECT  18.34 385.14 18.9 385.98 ;
     RECT  604.66 385.42 605.78 385.98 ;
     RECT  18.62 385.98 18.9 386.26 ;
     RECT  605.5 385.98 605.78 386.26 ;
     RECT  95 385.42 531.39 600.88 ;
     RECT  31.41 382.62 38.59 605.374 ;
     RECT  76.21 380.38 83.39 605.374 ;
     RECT  121.01 600.88 128.19 605.374 ;
     RECT  165.81 600.88 172.99 605.374 ;
     RECT  210.61 600.88 217.79 605.374 ;
     RECT  255.41 600.88 262.59 605.374 ;
     RECT  300.21 600.88 307.39 605.374 ;
     RECT  345.01 600.88 352.19 605.374 ;
     RECT  389.81 600.88 396.99 605.374 ;
     RECT  434.61 600.88 441.79 605.374 ;
     RECT  479.41 600.88 486.59 605.374 ;
     RECT  524.21 600.88 531.39 605.374 ;
     RECT  569.01 370.86 576.19 605.374 ;
     RECT  36.45 605.374 38.59 610.414 ;
     RECT  81.25 605.374 83.39 610.414 ;
     RECT  126.05 605.374 128.19 610.414 ;
     RECT  170.85 605.374 172.99 610.414 ;
     RECT  215.65 605.374 217.79 610.414 ;
     RECT  260.45 605.374 262.59 610.414 ;
     RECT  305.25 605.374 307.39 610.414 ;
     RECT  350.05 605.374 352.19 610.414 ;
     RECT  394.85 605.374 396.99 610.414 ;
     RECT  439.65 605.374 441.79 610.414 ;
     RECT  484.45 605.374 486.59 610.414 ;
     RECT  529.25 605.374 531.39 610.414 ;
     RECT  574.05 605.374 576.19 610.414 ;
    LAYER Metal3 ;
     RECT  0.26 364.42 13.02 372.54 ;
     RECT  13.02 364.42 13.3 382.62 ;
     RECT  13.3 365.54 18.06 382.62 ;
     RECT  18.06 367.78 31.954 382.62 ;
     RECT  31.954 9.556 32.926 605.324 ;
     RECT  32.926 14.596 37.074 605.324 ;
     RECT  37.074 14.596 38.246 610.364 ;
     RECT  58.66 356.58 76.834 356.86 ;
     RECT  76.834 9.556 77.846 605.324 ;
     RECT  77.846 14.596 81.454 605.324 ;
     RECT  81.454 14.596 82.766 610.364 ;
     RECT  82.766 14.596 90.02 19.18 ;
     RECT  90.02 13.3 95 19.18 ;
     RECT  82.766 218.26 95 220.78 ;
     RECT  82.766 260.26 95 260.54 ;
     RECT  82.766 348.74 95 356.86 ;
     RECT  95 13.3 100.94 260.54 ;
     RECT  100.94 9.38 112.36 260.54 ;
     RECT  112.36 8.26 112.83 260.54 ;
     RECT  112.83 9.556 121.634 260.54 ;
     RECT  95 348.74 121.634 600.88 ;
     RECT  121.634 9.556 122.846 605.324 ;
     RECT  122.846 13.3 126.454 605.324 ;
     RECT  126.454 13.3 127.566 610.364 ;
     RECT  127.566 13.3 144.34 252.88 ;
     RECT  144.34 12.74 147.98 252.88 ;
     RECT  147.98 11.62 157.5 252.88 ;
     RECT  157.5 9.38 166.054 252.88 ;
     RECT  127.566 348.74 166.054 349.58 ;
     RECT  127.566 368 166.054 600.88 ;
     RECT  166.054 9.38 166.36 605.324 ;
     RECT  166.36 8.26 168.14 605.324 ;
     RECT  168.14 13.3 171.454 605.324 ;
     RECT  171.454 13.3 172.366 610.364 ;
     RECT  172.366 13.3 205.77 252.88 ;
     RECT  205.77 6.58 206.24 252.88 ;
     RECT  172.366 348.74 207.62 349.58 ;
     RECT  206.24 9.38 211.054 252.88 ;
     RECT  207.62 348.74 211.054 351.26 ;
     RECT  172.366 368 211.054 600.88 ;
     RECT  211.054 9.38 216.02 605.324 ;
     RECT  216.02 13.3 216.274 605.324 ;
     RECT  216.274 13.3 217.346 610.364 ;
     RECT  217.346 348.74 235.34 351.26 ;
     RECT  217.346 13.3 251.67 252.88 ;
     RECT  251.67 8.82 256.034 252.88 ;
     RECT  235.34 348.74 256.034 349.58 ;
     RECT  217.346 368 256.034 600.88 ;
     RECT  256.034 8.82 258.16 605.324 ;
     RECT  258.16 8.26 259.42 605.324 ;
     RECT  259.42 12.18 261.074 605.324 ;
     RECT  261.074 12.18 262.346 610.364 ;
     RECT  262.346 12.18 268.38 252.88 ;
     RECT  268.38 16.1 297.76 252.88 ;
     RECT  297.76 9.38 298.9 252.88 ;
     RECT  298.9 9.556 300.834 252.88 ;
     RECT  262.346 348.74 300.834 349.02 ;
     RECT  262.346 368 300.834 600.88 ;
     RECT  300.834 9.556 301.946 605.324 ;
     RECT  301.946 14.596 305.554 605.324 ;
     RECT  305.554 14.596 306.766 610.364 ;
     RECT  306.766 20 345.634 252.88 ;
     RECT  306.766 368 345.634 600.88 ;
     RECT  345.634 9.556 346.946 605.324 ;
     RECT  346.946 13.3 350.554 605.324 ;
     RECT  350.554 13.3 351.566 610.364 ;
     RECT  351.566 13.3 360.76 252.88 ;
     RECT  360.76 8.82 361.62 252.88 ;
     RECT  351.566 348.74 367.78 349.02 ;
     RECT  367.78 348.74 371.14 349.58 ;
     RECT  371.14 348.74 376.74 350.7 ;
     RECT  361.62 12.18 377.67 252.88 ;
     RECT  377.67 8.82 378 252.88 ;
     RECT  378 12.18 390.154 252.88 ;
     RECT  376.74 348.74 390.154 351.26 ;
     RECT  351.566 368 390.154 600.88 ;
     RECT  390.154 9.556 395.474 605.324 ;
     RECT  395.474 9.556 396.446 610.364 ;
     RECT  396.446 9.556 399.98 252.88 ;
     RECT  399.98 9.38 409.36 252.88 ;
     RECT  409.36 8.82 410.06 252.88 ;
     RECT  396.446 348.74 411.74 351.26 ;
     RECT  410.06 13.3 435.154 252.88 ;
     RECT  411.74 348.74 435.154 349.58 ;
     RECT  396.446 368 435.154 600.88 ;
     RECT  435.154 9.556 436.126 605.324 ;
     RECT  436.126 11.62 440.274 605.324 ;
     RECT  440.274 11.62 441.446 610.364 ;
     RECT  441.446 11.62 450.76 252.88 ;
     RECT  450.76 8.26 457.1 252.88 ;
     RECT  457.1 9.38 461.3 252.88 ;
     RECT  441.446 348.74 470.26 349.58 ;
     RECT  461.3 11.62 480.034 252.88 ;
     RECT  470.26 348.74 480.034 356.3 ;
     RECT  441.446 368 480.034 600.88 ;
     RECT  480.034 9.556 481.046 605.324 ;
     RECT  481.046 12.74 484.654 605.324 ;
     RECT  484.654 12.74 485.66 610.364 ;
     RECT  485.66 13.3 485.966 610.364 ;
     RECT  485.966 348.74 499.38 356.3 ;
     RECT  485.966 368 499.38 600.88 ;
     RECT  499.38 348.74 510.3 600.88 ;
     RECT  485.966 13.3 511.96 252.88 ;
     RECT  511.96 11.62 524.834 252.88 ;
     RECT  510.3 348.74 524.834 356.3 ;
     RECT  510.3 368 524.834 600.88 ;
     RECT  524.834 9.556 526.046 605.324 ;
     RECT  526.046 13.3 529.654 605.324 ;
     RECT  529.654 13.3 530.766 610.364 ;
     RECT  530.766 348.74 532.14 349.58 ;
     RECT  530.766 13.3 537.74 13.58 ;
     RECT  532.14 348.74 537.74 349.02 ;
     RECT  569.254 9.556 570.526 605.324 ;
     RECT  570.526 14.596 574.654 605.324 ;
     RECT  574.654 14.596 575.566 610.364 ;
     RECT  590.38 372.82 596.26 373.1 ;
     RECT  596.26 369.46 599.9 373.1 ;
     RECT  599.9 363.3 604.1 373.1 ;
     RECT  604.1 363.3 606.06 378.14 ;
     RECT  606.06 363.3 613.04 373.66 ;
     RECT  613.04 363.3 615.58 372.54 ;
     RECT  615.58 364.42 619.74 372.54 ;
    LAYER Metal4 ;
     RECT  159.98 0.9 162.22 1.12 ;
     RECT  249.98 0.9 252.22 1.12 ;
     RECT  372.38 0.9 376.42 1.12 ;
     RECT  505.58 0.9 510.52 1.12 ;
     RECT  504.68 1.12 512.32 1.9 ;
     RECT  205.88 1.12 215.32 6.94 ;
     RECT  360.68 1.12 377.32 8.74 ;
     RECT  234.68 1.12 267.52 9.18 ;
     RECT  402.08 1.12 409.72 9.18 ;
     RECT  105.08 1.12 112.72 9.506 ;
     RECT  153.68 1.12 166.72 9.506 ;
     RECT  297.68 1.12 298.12 9.506 ;
     RECT  360.68 8.74 378.22 9.506 ;
     RECT  402.08 9.18 402.52 9.506 ;
     RECT  450.68 1.12 463.72 9.506 ;
     RECT  510.08 1.9 512.32 9.506 ;
     RECT  105.08 9.506 124.32 9.74 ;
     RECT  297.68 9.506 303.52 9.74 ;
     RECT  343.84 9.506 402.52 9.74 ;
     RECT  433.44 9.506 482.72 11.98 ;
     RECT  254.24 9.18 267.52 12.54 ;
     RECT  343.84 9.74 398.16 12.54 ;
     RECT  463.28 11.98 482.72 12.54 ;
     RECT  153.68 9.506 169.12 13.1 ;
     RECT  510.08 9.506 527.52 13.1 ;
     RECT  30.24 9.506 34.72 14.546 ;
     RECT  75.04 9.506 79.52 14.546 ;
     RECT  119.84 9.74 124.32 14.546 ;
     RECT  164.64 13.1 169.12 14.546 ;
     RECT  209.44 6.94 215.32 14.546 ;
     RECT  234.68 9.18 235.12 14.546 ;
     RECT  299.04 9.74 303.52 14.546 ;
     RECT  478.24 12.54 482.72 14.546 ;
     RECT  523.04 13.1 527.52 14.546 ;
     RECT  567.84 9.506 572.32 14.546 ;
     RECT  209.44 14.546 235.12 19.26 ;
     RECT  30.24 14.546 39.76 605.374 ;
     RECT  75.04 14.546 84.56 605.374 ;
     RECT  119.84 14.546 129.36 605.374 ;
     RECT  164.64 14.546 174.16 605.374 ;
     RECT  209.44 19.26 218.96 605.374 ;
     RECT  254.24 12.54 263.76 605.374 ;
     RECT  299.04 14.546 308.56 605.374 ;
     RECT  343.84 12.54 353.36 605.374 ;
     RECT  388.64 12.54 398.16 605.374 ;
     RECT  433.44 11.98 442.96 605.374 ;
     RECT  478.24 14.546 487.76 605.374 ;
     RECT  523.04 14.546 532.56 605.374 ;
     RECT  567.84 14.546 577.36 605.374 ;
     RECT  35.28 605.374 39.76 610.414 ;
     RECT  80.08 605.374 84.56 610.414 ;
     RECT  124.88 605.374 129.36 610.414 ;
     RECT  169.68 605.374 174.16 610.414 ;
     RECT  214.48 605.374 218.96 610.414 ;
     RECT  259.28 605.374 263.76 610.414 ;
     RECT  304.08 605.374 308.56 610.414 ;
     RECT  348.88 605.374 353.36 610.414 ;
     RECT  393.68 605.374 398.16 610.414 ;
     RECT  438.48 605.374 442.96 610.414 ;
     RECT  483.28 605.374 487.76 610.414 ;
     RECT  528.08 605.374 532.56 610.414 ;
     RECT  572.88 605.374 577.36 610.414 ;
  END
END mem_64_16_gf180
END LIBRARY
